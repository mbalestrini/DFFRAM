* NGSPICE file created from DFFRF_2R1W.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_2 abstract view
.subckt sky130_fd_sc_hd__ebufn_2 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlclkp_1 abstract view
.subckt sky130_fd_sc_hd__dlclkp_1 CLK GATE VGND VNB VPB VPWR GCLK
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_2 abstract view
.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

.subckt DFFRF_2R1W CLK DA[0] DA[10] DA[11] DA[12] DA[13] DA[14] DA[15] DA[16] DA[17]
+ DA[18] DA[19] DA[1] DA[20] DA[21] DA[22] DA[23] DA[24] DA[25] DA[26] DA[27] DA[28]
+ DA[29] DA[2] DA[30] DA[31] DA[3] DA[4] DA[5] DA[6] DA[7] DA[8] DA[9] DB[0] DB[10]
+ DB[11] DB[12] DB[13] DB[14] DB[15] DB[16] DB[17] DB[18] DB[19] DB[1] DB[20] DB[21]
+ DB[22] DB[23] DB[24] DB[25] DB[26] DB[27] DB[28] DB[29] DB[2] DB[30] DB[31] DB[3]
+ DB[4] DB[5] DB[6] DB[7] DB[8] DB[9] DW[0] DW[10] DW[11] DW[12] DW[13] DW[14] DW[15]
+ DW[16] DW[17] DW[18] DW[19] DW[1] DW[20] DW[21] DW[22] DW[23] DW[24] DW[25] DW[26]
+ DW[27] DW[28] DW[29] DW[2] DW[30] DW[31] DW[3] DW[4] DW[5] DW[6] DW[7] DW[8] DW[9]
+ RA[0] RA[1] RA[2] RA[3] RA[4] RB[0] RB[1] RB[2] RB[3] RB[4] RW[0] RW[1] RW[2] RW[3]
+ RW[4] VGND VPWR WE
Xtap_24_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_40_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[21\].RFW.BIT\[12\].FF REGF\[21\].RFW.CG\[1\]/GCLK DW[12] VGND VGND VPWR VPWR
+ REGF\[21\].RFW.BIT\[12\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_12_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_12_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_12_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[10\].RFW.BIT\[13\].OBUF2 REGF\[10\].RFW.BIT\[13\].FF/Q REGF\[10\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[13] sky130_fd_sc_hd__ebufn_2
Xtap_22_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_37_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_37_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_37_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_37_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_37_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[8\].RFW.BIT\[28\].OBUF1 REGF\[8\].RFW.BIT\[28\].FF/Q REGF\[8\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[28] sky130_fd_sc_hd__ebufn_2
XREGF\[10\].RFW.BIT\[25\].FF REGF\[10\].RFW.CG\[3\]/GCLK DW[25] VGND VGND VPWR VPWR
+ REGF\[10\].RFW.BIT\[25\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_53_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_53_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_53_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_53_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_9_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_9_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_9_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDEC2.D.AND2 RW[3] RW[4] DEC2.TIE/HI VGND VGND VPWR VPWR DEC2.D.AND2/X sky130_fd_sc_hd__and3b_4
XREGF\[26\].RFW.BIT\[23\].OBUF1 REGF\[26\].RFW.BIT\[23\].FF/Q REGF\[26\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[23] sky130_fd_sc_hd__ebufn_2
Xfill_9_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_9_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[31\].RFW.BIT\[12\].OBUF1 REGF\[31\].RFW.BIT\[12\].FF/Q REGF\[31\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[12] sky130_fd_sc_hd__ebufn_2
Xfill_50_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_43_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_36_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[21\].RFW.BIT\[1\].FF REGF\[21\].RFW.CG\[0\]/GCLK DW[1] VGND VGND VPWR VPWR
+ REGF\[21\].RFW.BIT\[1\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_29_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_58_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_58_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[3\].FF REGF\[20\].RFW.CG\[0\]/GCLK DW[3] VGND VGND VPWR VPWR
+ REGF\[20\].RFW.BIT\[3\].FF/Q sky130_fd_sc_hd__dfxtp_1
XDEC0.D0.ABUF\[2\] RA[2] VGND VGND VPWR VPWR DEC0.D0.AND7/C sky130_fd_sc_hd__clkbuf_2
XREGF\[22\].RFW.BIT\[26\].OBUF1 REGF\[22\].RFW.BIT\[26\].FF/Q REGF\[22\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[26] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.CG\[2\] CLK REGF\[26\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[26\].RFW.CG\[2\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_1_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[7\].RFW.BIT\[16\].OBUF1 REGF\[7\].RFW.BIT\[16\].FF/Q REGF\[7\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[16] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[18\].FF REGF\[5\].RFW.CG\[2\]/GCLK DW[18] VGND VGND VPWR VPWR
+ REGF\[5\].RFW.BIT\[18\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[1\].RFW.BIT\[20\].FF REGF\[1\].RFW.CG\[2\]/GCLK DW[20] VGND VGND VPWR VPWR
+ REGF\[1\].RFW.BIT\[20\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_23_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_23_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_23_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_23_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[25\].RFW.BIT\[11\].OBUF1 REGF\[25\].RFW.BIT\[11\].FF/Q REGF\[25\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[11] sky130_fd_sc_hd__ebufn_2
Xfill_48_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_48_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[7\].RFW.INV2\[3\] DEC1.D0.AND7/X VGND VGND VPWR VPWR REGF\[7\].RFW.INV2\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[5\].RFW.BIT\[0\].FF REGF\[5\].RFW.CG\[0\]/GCLK DW[0] VGND VGND VPWR VPWR REGF\[5\].RFW.BIT\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[26\].RFW.BIT\[27\].OBUF2 REGF\[26\].RFW.BIT\[27\].FF/Q REGF\[26\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[27] sky130_fd_sc_hd__ebufn_2
Xfill_22_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_15_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[31\].RFW.BIT\[16\].OBUF2 REGF\[31\].RFW.BIT\[16\].FF/Q REGF\[31\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[16] sky130_fd_sc_hd__ebufn_2
XREGF\[31\].RFW.BIT\[0\].OBUF1 REGF\[31\].RFW.BIT\[0\].FF/Q REGF\[31\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[0] sky130_fd_sc_hd__ebufn_2
XREGF\[22\].RFW.BIT\[18\].FF REGF\[22\].RFW.CG\[2\]/GCLK DW[18] VGND VGND VPWR VPWR
+ REGF\[22\].RFW.BIT\[18\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[3\].RFW.BIT\[19\].OBUF1 REGF\[3\].RFW.BIT\[19\].FF/Q REGF\[3\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[19] sky130_fd_sc_hd__ebufn_2
XREGF\[11\].RFW.INV2\[0\] DEC1.D1.AND3/X VGND VGND VPWR VPWR REGF\[11\].RFW.INV2\[0\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[28\].RFW.BIT\[12\].FF REGF\[28\].RFW.CG\[1\]/GCLK DW[12] VGND VGND VPWR VPWR
+ REGF\[28\].RFW.BIT\[12\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[16\].RFW.BIT\[25\].OBUF1 REGF\[16\].RFW.BIT\[25\].FF/Q REGF\[16\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[25] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.BIT\[12\].OBUF2 REGF\[29\].RFW.BIT\[12\].FF/Q REGF\[29\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[12] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.INV2\[1\] DEC1.D3.AND3/X VGND VGND VPWR VPWR REGF\[27\].RFW.INV2\[1\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[4\].RFW.BIT\[2\].FF REGF\[4\].RFW.CG\[0\]/GCLK DW[2] VGND VGND VPWR VPWR REGF\[4\].RFW.BIT\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[21\].RFW.BIT\[14\].OBUF1 REGF\[21\].RFW.BIT\[14\].FF/Q REGF\[21\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[14] sky130_fd_sc_hd__ebufn_2
Xfill_41_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[19\].RFW.BIT\[10\].OBUF1 REGF\[19\].RFW.BIT\[10\].FF/Q REGF\[19\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[10] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.BIT\[25\].FF REGF\[17\].RFW.CG\[3\]/GCLK DW[25] VGND VGND VPWR VPWR
+ REGF\[17\].RFW.BIT\[25\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[14\].RFW.CG\[2\] CLK REGF\[14\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[14\].RFW.CG\[2\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[3\].RFW.BIT\[4\].FF REGF\[3\].RFW.CG\[0\]/GCLK DW[4] VGND VGND VPWR VPWR REGF\[3\].RFW.BIT\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xtap_56_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_46_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.BIT\[28\].OBUF1 REGF\[12\].RFW.BIT\[28\].FF/Q REGF\[12\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[28] sky130_fd_sc_hd__ebufn_2
Xfill_18_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[25\].RFW.BIT\[15\].OBUF2 REGF\[25\].RFW.BIT\[15\].FF/Q REGF\[25\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[15] sky130_fd_sc_hd__ebufn_2
Xfill_18_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_18_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_62_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[2\].RFW.BIT\[6\].FF REGF\[2\].RFW.CG\[0\]/GCLK DW[6] VGND VGND VPWR VPWR REGF\[2\].RFW.BIT\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[31\].RFW.BIT\[7\].FF REGF\[31\].RFW.CG\[0\]/GCLK DW[7] VGND VGND VPWR VPWR
+ REGF\[31\].RFW.BIT\[7\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_34_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.BIT\[20\].OBUF1 REGF\[3\].RFW.BIT\[20\].FF/Q REGF\[3\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[20] sky130_fd_sc_hd__ebufn_2
XREGF\[23\].RFW.INV1\[2\] DEC0.D2.AND7/X VGND VGND VPWR VPWR REGF\[23\].RFW.INV1\[2\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_50_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_50_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[15\].RFW.BIT\[13\].OBUF1 REGF\[15\].RFW.BIT\[13\].FF/Q REGF\[15\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[13] sky130_fd_sc_hd__ebufn_2
Xfill_6_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[30\].RFW.BIT\[9\].FF REGF\[30\].RFW.CG\[1\]/GCLK DW[9] VGND VGND VPWR VPWR
+ REGF\[30\].RFW.BIT\[9\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_59_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_59_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_59_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_6_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_6_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[1\].RFW.BIT\[8\].FF REGF\[1\].RFW.CG\[1\]/GCLK DW[8] VGND VGND VPWR VPWR REGF\[1\].RFW.BIT\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[31\].RFW.BIT\[4\].OBUF2 REGF\[31\].RFW.BIT\[4\].FF/Q REGF\[31\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[4] sky130_fd_sc_hd__ebufn_2
Xgenblk1.RFW0.BIT\[29\].OBUF1 genblk1.RFW0.TIE\[3\]/LO genblk1.RFW0.INV1\[3\]/Y VGND
+ VGND VPWR VPWR DA[29] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[29\].OBUF2 REGF\[16\].RFW.BIT\[29\].FF/Q REGF\[16\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[29] sky130_fd_sc_hd__ebufn_2
Xfill_20_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_13_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[2\].RFW.BIT\[26\].FF REGF\[2\].RFW.CG\[3\]/GCLK DW[26] VGND VGND VPWR VPWR
+ REGF\[2\].RFW.BIT\[26\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[21\].RFW.BIT\[18\].OBUF2 REGF\[21\].RFW.BIT\[18\].FF/Q REGF\[21\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[18] sky130_fd_sc_hd__ebufn_2
XREGF\[22\].RFW.BIT\[31\].OBUF2 REGF\[22\].RFW.BIT\[31\].FF/Q REGF\[22\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[31] sky130_fd_sc_hd__ebufn_2
XREGF\[8\].RFW.BIT\[20\].FF REGF\[8\].RFW.CG\[2\]/GCLK DW[20] VGND VGND VPWR VPWR
+ REGF\[8\].RFW.BIT\[20\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[7\].RFW.BIT\[21\].OBUF2 REGF\[7\].RFW.BIT\[21\].FF/Q REGF\[7\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[21] sky130_fd_sc_hd__ebufn_2
XREGF\[14\].RFW.BIT\[10\].FF REGF\[14\].RFW.CG\[1\]/GCLK DW[10] VGND VGND VPWR VPWR
+ REGF\[14\].RFW.BIT\[10\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[30\].RFW.BIT\[13\].FF REGF\[30\].RFW.CG\[1\]/GCLK DW[13] VGND VGND VPWR VPWR
+ REGF\[30\].RFW.BIT\[13\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[19\].RFW.BIT\[14\].OBUF2 REGF\[19\].RFW.BIT\[14\].FF/Q REGF\[19\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[14] sky130_fd_sc_hd__ebufn_2
XREGF\[11\].RFW.BIT\[16\].OBUF1 REGF\[11\].RFW.BIT\[16\].FF/Q REGF\[11\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[16] sky130_fd_sc_hd__ebufn_2
XDEC2.D2.ABUF\[0\] RW[0] VGND VGND VPWR VPWR DEC2.D2.AND7/A sky130_fd_sc_hd__clkbuf_2
XREGF\[29\].RFW.BIT\[18\].FF REGF\[29\].RFW.CG\[2\]/GCLK DW[18] VGND VGND VPWR VPWR
+ REGF\[29\].RFW.BIT\[18\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_54_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[25\].RFW.BIT\[20\].FF REGF\[25\].RFW.CG\[2\]/GCLK DW[20] VGND VGND VPWR VPWR
+ REGF\[25\].RFW.BIT\[20\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_20_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_20_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_20_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_47_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_29_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_29_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgenblk1.RFW0.BIT\[30\].OBUF1 genblk1.RFW0.TIE\[3\]/LO genblk1.RFW0.INV1\[3\]/Y VGND
+ VGND VPWR VPWR DA[30] sky130_fd_sc_hd__ebufn_2
Xfill_29_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_29_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_29_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.BIT\[24\].OBUF2 REGF\[3\].RFW.BIT\[24\].FF/Q REGF\[3\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[24] sky130_fd_sc_hd__ebufn_2
XREGF\[15\].RFW.BIT\[17\].OBUF2 REGF\[15\].RFW.BIT\[17\].FF/Q REGF\[15\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[17] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[30\].OBUF2 REGF\[16\].RFW.BIT\[30\].FF/Q REGF\[16\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[30] sky130_fd_sc_hd__ebufn_2
Xfill_45_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_45_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_45_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_45_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_45_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.INV1\[3\] DEC0.D2.AND2/X VGND VGND VPWR VPWR REGF\[18\].RFW.INV1\[3\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_61_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_61_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_61_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_61_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xgenblk1.RFW0.TIE\[4\] VGND VGND VPWR VPWR genblk1.RFW0.TIE\[4\]/HI genblk1.RFW0.TIE\[4\]/LO
+ sky130_fd_sc_hd__conb_1
Xfill_11_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_9_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_40_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[2\].RFW.BIT\[12\].OBUF2 REGF\[2\].RFW.BIT\[12\].FF/Q REGF\[2\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[12] sky130_fd_sc_hd__ebufn_2
Xfill_15_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_15_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XREGF\[22\].RFW.CGAND DEC2.D2.AND6/X WE VGND VGND VPWR VPWR REGF\[22\].RFW.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_15_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_15_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_15_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[9\].RFW.BIT\[26\].FF REGF\[9\].RFW.CG\[3\]/GCLK DW[26] VGND VGND VPWR VPWR
+ REGF\[9\].RFW.BIT\[26\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[15\].RFW.BIT\[16\].FF REGF\[15\].RFW.CG\[2\]/GCLK DW[16] VGND VGND VPWR VPWR
+ REGF\[15\].RFW.BIT\[16\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_31_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_52_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_31_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_31_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_31_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.BIT\[19\].FF REGF\[31\].RFW.CG\[2\]/GCLK DW[19] VGND VGND VPWR VPWR
+ REGF\[31\].RFW.BIT\[19\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[9\].RFW.INV2\[0\] DEC1.D1.AND1/X VGND VGND VPWR VPWR REGF\[9\].RFW.INV2\[0\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_56_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_56_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_3_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_3_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[11\].RFW.BIT\[21\].OBUF2 REGF\[11\].RFW.BIT\[21\].FF/Q REGF\[11\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[21] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[26\].FF REGF\[26\].RFW.CG\[3\]/GCLK DW[26] VGND VGND VPWR VPWR
+ REGF\[26\].RFW.BIT\[26\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[30\].RFW.BIT\[2\].OBUF2 REGF\[30\].RFW.BIT\[2\].FF/Q REGF\[30\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[2] sky130_fd_sc_hd__ebufn_2
Xfill_59_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[26\].RFW.BIT\[18\].OBUF1 REGF\[26\].RFW.BIT\[18\].FF/Q REGF\[26\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[18] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[31\].OBUF1 REGF\[27\].RFW.BIT\[31\].FF/Q REGF\[27\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[31] sky130_fd_sc_hd__ebufn_2
Xfill_7_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[5\].RFW.INV1\[1\] DEC0.D0.AND5/X VGND VGND VPWR VPWR REGF\[5\].RFW.INV1\[1\]/Y
+ sky130_fd_sc_hd__inv_4
XDEC1.D3.ABUF\[1\] RB[1] VGND VGND VPWR VPWR DEC1.D3.AND7/B sky130_fd_sc_hd__clkbuf_2
XREGF\[6\].RFW.BIT\[11\].FF REGF\[6\].RFW.CG\[1\]/GCLK DW[11] VGND VGND VPWR VPWR
+ REGF\[6\].RFW.BIT\[11\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_31_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_38_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_54_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_26_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_26_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_26_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_42_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_42_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_42_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[8\].RFW.BIT\[24\].OBUF1 REGF\[8\].RFW.BIT\[24\].FF/Q REGF\[8\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[24] sky130_fd_sc_hd__ebufn_2
XREGF\[23\].RFW.BIT\[11\].FF REGF\[23\].RFW.CG\[1\]/GCLK DW[11] VGND VGND VPWR VPWR
+ REGF\[23\].RFW.BIT\[11\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_52_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_45_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_38_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_0_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC2.D1.AND7 DEC2.D1.AND7/A DEC2.D1.AND7/B DEC2.D1.AND7/C DEC2.D1.AND7/D VGND VGND
+ VPWR VPWR DEC2.D1.AND7/X sky130_fd_sc_hd__and4_2
XREGF\[12\].RFW.BIT\[24\].FF REGF\[12\].RFW.CG\[3\]/GCLK DW[24] VGND VGND VPWR VPWR
+ REGF\[12\].RFW.BIT\[24\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[22\].RFW.CG\[1\] CLK REGF\[22\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[22\].RFW.CG\[1\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[4\].RFW.BIT\[27\].OBUF1 REGF\[4\].RFW.BIT\[27\].FF/Q REGF\[4\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[27] sky130_fd_sc_hd__ebufn_2
XREGF\[22\].RFW.BIT\[22\].OBUF1 REGF\[22\].RFW.BIT\[22\].FF/Q REGF\[22\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[22] sky130_fd_sc_hd__ebufn_2
Xfill_12_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_12_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_12_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[7\].RFW.BIT\[12\].OBUF1 REGF\[7\].RFW.BIT\[12\].FF/Q REGF\[7\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[12] sky130_fd_sc_hd__ebufn_2
Xtap_22_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_37_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_37_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_37_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_37_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_37_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_37_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[8\].RFW.BIT\[28\].OBUF2 REGF\[8\].RFW.BIT\[28\].FF/Q REGF\[8\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[28] sky130_fd_sc_hd__ebufn_2
Xfill_53_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_53_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_53_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_53_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_53_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_9_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_9_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC2.D.AND3 RW[4] RW[3] DEC2.TIE/HI VGND VGND VPWR VPWR DEC2.D.AND3/X sky130_fd_sc_hd__and3_4
XREGF\[26\].RFW.BIT\[23\].OBUF2 REGF\[26\].RFW.BIT\[23\].FF/Q REGF\[26\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[23] sky130_fd_sc_hd__ebufn_2
Xfill_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_9_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_9_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[7\].RFW.BIT\[17\].FF REGF\[7\].RFW.CG\[2\]/GCLK DW[17] VGND VGND VPWR VPWR
+ REGF\[7\].RFW.BIT\[17\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[31\].RFW.BIT\[12\].OBUF2 REGF\[31\].RFW.BIT\[12\].FF/Q REGF\[31\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[12] sky130_fd_sc_hd__ebufn_2
Xfill_50_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_43_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.BIT\[15\].OBUF1 REGF\[3\].RFW.BIT\[15\].FF/Q REGF\[3\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[15] sky130_fd_sc_hd__ebufn_2
Xfill_36_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[16\].RFW.BIT\[21\].OBUF1 REGF\[16\].RFW.BIT\[21\].FF/Q REGF\[16\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[21] sky130_fd_sc_hd__ebufn_2
Xfill_29_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XREGF\[10\].RFW.CG\[1\] CLK REGF\[10\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[10\].RFW.CG\[1\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[21\].RFW.BIT\[10\].OBUF1 REGF\[21\].RFW.BIT\[10\].FF/Q REGF\[21\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[10] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[17\].FF REGF\[24\].RFW.CG\[2\]/GCLK DW[17] VGND VGND VPWR VPWR
+ REGF\[24\].RFW.BIT\[17\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[22\].RFW.BIT\[26\].OBUF2 REGF\[22\].RFW.BIT\[26\].FF/Q REGF\[22\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[26] sky130_fd_sc_hd__ebufn_2
XREGF\[7\].RFW.BIT\[16\].OBUF2 REGF\[7\].RFW.BIT\[16\].FF/Q REGF\[7\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[16] sky130_fd_sc_hd__ebufn_2
XREGF\[31\].RFW.INV1\[2\] DEC0.D3.AND7/X VGND VGND VPWR VPWR REGF\[31\].RFW.INV1\[2\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_23_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_23_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_23_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_23_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_23_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.BIT\[24\].OBUF1 REGF\[12\].RFW.BIT\[24\].FF/Q REGF\[12\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[24] sky130_fd_sc_hd__ebufn_2
XREGF\[25\].RFW.BIT\[11\].OBUF2 REGF\[25\].RFW.BIT\[11\].FF/Q REGF\[25\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[11] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.BIT\[24\].FF REGF\[19\].RFW.CG\[3\]/GCLK DW[24] VGND VGND VPWR VPWR
+ REGF\[19\].RFW.BIT\[24\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_48_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_48_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[14\].RFW.INV2\[1\] DEC1.D1.AND6/X VGND VGND VPWR VPWR REGF\[14\].RFW.INV2\[1\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_22_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_15_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.BIT\[0\].OBUF2 REGF\[31\].RFW.BIT\[0\].FF/Q REGF\[31\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[0] sky130_fd_sc_hd__ebufn_2
Xgenblk1.RFW0.BIT\[25\].OBUF1 genblk1.RFW0.TIE\[3\]/LO genblk1.RFW0.INV1\[3\]/Y VGND
+ VGND VPWR VPWR DA[25] sky130_fd_sc_hd__ebufn_2
XREGF\[3\].RFW.BIT\[19\].OBUF2 REGF\[3\].RFW.BIT\[19\].FF/Q REGF\[3\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[19] sky130_fd_sc_hd__ebufn_2
XDEC0.D2.AND0 DEC0.D2.AND7/A DEC0.D2.AND7/B DEC0.D2.AND7/C DEC0.D2.AND7/D VGND VGND
+ VPWR VPWR DEC0.D2.AND0/Y sky130_fd_sc_hd__nor4b_2
XREGF\[16\].RFW.BIT\[25\].OBUF2 REGF\[16\].RFW.BIT\[25\].FF/Q REGF\[16\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[25] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.BIT\[14\].OBUF2 REGF\[21\].RFW.BIT\[14\].FF/Q REGF\[21\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[14] sky130_fd_sc_hd__ebufn_2
Xfill_41_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_34_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[19\].RFW.BIT\[10\].OBUF2 REGF\[19\].RFW.BIT\[10\].FF/Q REGF\[19\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[10] sky130_fd_sc_hd__ebufn_2
XREGF\[11\].RFW.BIT\[12\].OBUF1 REGF\[11\].RFW.BIT\[12\].FF/Q REGF\[11\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[12] sky130_fd_sc_hd__ebufn_2
Xtap_56_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[10\].RFW.BIT\[15\].FF REGF\[10\].RFW.CG\[1\]/GCLK DW[15] VGND VGND VPWR VPWR
+ REGF\[10\].RFW.BIT\[15\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[4\].RFW.BIT\[25\].FF REGF\[4\].RFW.CG\[3\]/GCLK DW[25] VGND VGND VPWR VPWR
+ REGF\[4\].RFW.BIT\[25\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[10\].RFW.INV1\[2\] DEC0.D1.AND2/X VGND VGND VPWR VPWR REGF\[10\].RFW.INV1\[2\]/Y
+ sky130_fd_sc_hd__inv_4
Xtap_46_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.BIT\[28\].OBUF2 REGF\[12\].RFW.BIT\[28\].FF/Q REGF\[12\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[28] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.INV1\[3\] DEC0.D3.AND2/X VGND VGND VPWR VPWR REGF\[26\].RFW.INV1\[3\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_18_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_18_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_18_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_62_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_34_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.BIT\[20\].OBUF2 REGF\[3\].RFW.BIT\[20\].FF/Q REGF\[3\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[20] sky130_fd_sc_hd__ebufn_2
Xfill_50_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_50_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_50_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[15\].RFW.BIT\[13\].OBUF2 REGF\[15\].RFW.BIT\[13\].FF/Q REGF\[15\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[13] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.BIT\[8\].FF REGF\[19\].RFW.CG\[1\]/GCLK DW[8] VGND VGND VPWR VPWR
+ REGF\[19\].RFW.BIT\[8\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_6_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[21\].RFW.BIT\[25\].FF REGF\[21\].RFW.CG\[3\]/GCLK DW[25] VGND VGND VPWR VPWR
+ REGF\[21\].RFW.BIT\[25\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_59_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_59_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_59_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_59_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_6_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_6_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgenblk1.RFW0.BIT\[29\].OBUF2 genblk1.RFW0.TIE\[7\]/LO genblk1.RFW0.INV2\[3\]/Y VGND
+ VGND VPWR VPWR DB[29] sky130_fd_sc_hd__ebufn_2
Xfill_20_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_13_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[11\].RFW.BIT\[16\].OBUF2 REGF\[11\].RFW.BIT\[16\].FF/Q REGF\[11\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[16] sky130_fd_sc_hd__ebufn_2
XREGF\[1\].RFW.BIT\[10\].FF REGF\[1\].RFW.CG\[1\]/GCLK DW[10] VGND VGND VPWR VPWR
+ REGF\[1\].RFW.BIT\[10\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[21\].RFW.CGAND DEC2.D2.AND5/X WE VGND VGND VPWR VPWR REGF\[21\].RFW.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xtap_54_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_20_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_20_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_20_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[27\].RFW.BIT\[26\].OBUF1 REGF\[27\].RFW.BIT\[26\].FF/Q REGF\[27\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[26] sky130_fd_sc_hd__ebufn_2
Xtap_47_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.CG\[3\] CLK REGF\[31\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[31\].RFW.CG\[3\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_29_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgenblk1.RFW0.BIT\[30\].OBUF2 genblk1.RFW0.TIE\[7\]/LO genblk1.RFW0.INV2\[3\]/Y VGND
+ VGND VPWR VPWR DB[30] sky130_fd_sc_hd__ebufn_2
Xfill_29_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_29_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_29_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_45_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_45_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_45_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_45_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_45_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_45_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_61_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_61_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_61_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_61_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_61_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[17\].RFW.BIT\[15\].FF REGF\[17\].RFW.CG\[1\]/GCLK DW[15] VGND VGND VPWR VPWR
+ REGF\[17\].RFW.BIT\[15\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[23\].RFW.BIT\[29\].OBUF1 REGF\[23\].RFW.BIT\[29\].FF/Q REGF\[23\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[29] sky130_fd_sc_hd__ebufn_2
XREGF\[30\].RFW.CG\[0\] CLK REGF\[30\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[30\].RFW.CG\[0\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_9_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[8\].RFW.BIT\[19\].OBUF1 REGF\[8\].RFW.BIT\[19\].FF/Q REGF\[8\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[19] sky130_fd_sc_hd__ebufn_2
Xfill_11_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XREGF\[26\].RFW.BIT\[14\].OBUF1 REGF\[26\].RFW.BIT\[14\].FF/Q REGF\[26\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[14] sky130_fd_sc_hd__ebufn_2
Xtap_26_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[28\].RFW.BIT\[25\].FF REGF\[28\].RFW.CG\[3\]/GCLK DW[25] VGND VGND VPWR VPWR
+ REGF\[28\].RFW.BIT\[25\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_15_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_15_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[8\].RFW.CG\[3\] CLK REGF\[8\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[8\].RFW.CG\[3\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_15_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_15_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_15_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_52_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_31_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_31_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_31_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_31_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_31_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_45_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[17\].RFW.BIT\[28\].OBUF1 REGF\[17\].RFW.BIT\[28\].FF/Q REGF\[17\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[28] sky130_fd_sc_hd__ebufn_2
XREGF\[2\].RFW.BIT\[16\].FF REGF\[2\].RFW.CG\[2\]/GCLK DW[16] VGND VGND VPWR VPWR
+ REGF\[2\].RFW.BIT\[16\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[22\].RFW.BIT\[17\].OBUF1 REGF\[22\].RFW.BIT\[17\].FF/Q REGF\[22\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[17] sky130_fd_sc_hd__ebufn_2
XREGF\[23\].RFW.BIT\[30\].OBUF1 REGF\[23\].RFW.BIT\[30\].FF/Q REGF\[23\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[30] sky130_fd_sc_hd__ebufn_2
Xfill_56_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_56_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_3_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[8\].RFW.BIT\[10\].FF REGF\[8\].RFW.CG\[1\]/GCLK DW[10] VGND VGND VPWR VPWR
+ REGF\[8\].RFW.BIT\[10\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_3_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[8\].RFW.BIT\[20\].OBUF1 REGF\[8\].RFW.BIT\[20\].FF/Q REGF\[8\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[20] sky130_fd_sc_hd__ebufn_2
XREGF\[7\].RFW.CG\[0\] CLK REGF\[7\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[7\].RFW.CG\[0\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[8\].RFW.INV1\[2\] DEC0.D1.AND0/Y VGND VGND VPWR VPWR REGF\[8\].RFW.INV1\[2\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_59_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[26\].RFW.BIT\[18\].OBUF2 REGF\[26\].RFW.BIT\[18\].FF/Q REGF\[26\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[18] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[31\].OBUF2 REGF\[27\].RFW.BIT\[31\].FF/Q REGF\[27\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[31] sky130_fd_sc_hd__ebufn_2
XREGF\[25\].RFW.BIT\[10\].FF REGF\[25\].RFW.CG\[1\]/GCLK DW[10] VGND VGND VPWR VPWR
+ REGF\[25\].RFW.BIT\[10\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_7_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[4\].RFW.BIT\[23\].OBUF1 REGF\[4\].RFW.BIT\[23\].FF/Q REGF\[4\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[23] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[16\].OBUF1 REGF\[16\].RFW.BIT\[16\].FF/Q REGF\[16\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[16] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.INV1\[0\] DEC0.D3.AND4/X VGND VGND VPWR VPWR REGF\[28\].RFW.INV1\[0\]/Y
+ sky130_fd_sc_hd__inv_4
Xtap_24_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[14\].RFW.BIT\[23\].FF REGF\[14\].RFW.CG\[2\]/GCLK DW[23] VGND VGND VPWR VPWR
+ REGF\[14\].RFW.BIT\[23\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_54_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[30\].RFW.BIT\[26\].FF REGF\[30\].RFW.CG\[3\]/GCLK DW[26] VGND VGND VPWR VPWR
+ REGF\[30\].RFW.BIT\[26\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_26_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_26_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_26_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_42_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_42_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_42_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[8\].RFW.BIT\[24\].OBUF2 REGF\[8\].RFW.BIT\[24\].FF/Q REGF\[8\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[24] sky130_fd_sc_hd__ebufn_2
Xfill_52_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.BIT\[19\].OBUF1 REGF\[12\].RFW.BIT\[19\].FF/Q REGF\[12\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[19] sky130_fd_sc_hd__ebufn_2
Xfill_45_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_38_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDEC1.D1.ABUF\[0\] RB[0] VGND VGND VPWR VPWR DEC1.D1.AND7/A sky130_fd_sc_hd__clkbuf_2
Xfill_0_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[16\].RFW.BIT\[1\].FF REGF\[16\].RFW.CG\[0\]/GCLK DW[1] VGND VGND VPWR VPWR
+ REGF\[16\].RFW.BIT\[1\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[3\].RFW.BIT\[11\].OBUF1 REGF\[3\].RFW.BIT\[11\].FF/Q REGF\[3\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[11] sky130_fd_sc_hd__ebufn_2
XREGF\[15\].RFW.BIT\[3\].FF REGF\[15\].RFW.CG\[0\]/GCLK DW[3] VGND VGND VPWR VPWR
+ REGF\[15\].RFW.BIT\[3\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[2\].RFW.INV2\[3\] DEC1.D0.AND2/X VGND VGND VPWR VPWR REGF\[2\].RFW.INV2\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[9\].RFW.BIT\[16\].FF REGF\[9\].RFW.CG\[2\]/GCLK DW[16] VGND VGND VPWR VPWR
+ REGF\[9\].RFW.BIT\[16\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[4\].RFW.BIT\[27\].OBUF2 REGF\[4\].RFW.BIT\[27\].FF/Q REGF\[4\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[27] sky130_fd_sc_hd__ebufn_2
XREGF\[22\].RFW.BIT\[22\].OBUF2 REGF\[22\].RFW.BIT\[22\].FF/Q REGF\[22\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[22] sky130_fd_sc_hd__ebufn_2
Xfill_12_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_12_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[14\].RFW.BIT\[5\].FF REGF\[14\].RFW.CG\[0\]/GCLK DW[5] VGND VGND VPWR VPWR
+ REGF\[14\].RFW.BIT\[5\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_12_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[7\].RFW.BIT\[12\].OBUF2 REGF\[7\].RFW.BIT\[12\].FF/Q REGF\[7\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[12] sky130_fd_sc_hd__ebufn_2
XREGF\[22\].RFW.INV2\[1\] DEC1.D2.AND6/X VGND VGND VPWR VPWR REGF\[22\].RFW.INV2\[1\]/Y
+ sky130_fd_sc_hd__inv_4
Xtap_22_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.BIT\[20\].OBUF1 REGF\[12\].RFW.BIT\[20\].FF/Q REGF\[12\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[20] sky130_fd_sc_hd__ebufn_2
Xfill_37_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_37_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_37_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[29\].RFW.BIT\[1\].FF REGF\[29\].RFW.CG\[0\]/GCLK DW[1] VGND VGND VPWR VPWR
+ REGF\[29\].RFW.BIT\[1\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_8_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[26\].RFW.BIT\[16\].FF REGF\[26\].RFW.CG\[2\]/GCLK DW[16] VGND VGND VPWR VPWR
+ REGF\[26\].RFW.BIT\[16\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_37_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_37_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_37_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_53_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_53_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[13\].RFW.BIT\[7\].FF REGF\[13\].RFW.CG\[0\]/GCLK DW[7] VGND VGND VPWR VPWR
+ REGF\[13\].RFW.BIT\[7\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_53_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_53_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_53_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_53_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_9_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_9_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_9_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_9_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_9_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[28\].RFW.BIT\[3\].FF REGF\[28\].RFW.CG\[0\]/GCLK DW[3] VGND VGND VPWR VPWR
+ REGF\[28\].RFW.BIT\[3\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[15\].RFW.BIT\[29\].FF REGF\[15\].RFW.CG\[3\]/GCLK DW[29] VGND VGND VPWR VPWR
+ REGF\[15\].RFW.BIT\[29\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_50_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[12\].RFW.BIT\[9\].FF REGF\[12\].RFW.CG\[1\]/GCLK DW[9] VGND VGND VPWR VPWR
+ REGF\[12\].RFW.BIT\[9\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[11\].RFW.BIT\[31\].FF REGF\[11\].RFW.CG\[3\]/GCLK DW[31] VGND VGND VPWR VPWR
+ REGF\[11\].RFW.BIT\[31\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xgenblk1.RFW0.BIT\[21\].OBUF1 genblk1.RFW0.TIE\[2\]/LO genblk1.RFW0.INV1\[2\]/Y VGND
+ VGND VPWR VPWR DA[21] sky130_fd_sc_hd__ebufn_2
Xfill_43_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[3\].RFW.BIT\[15\].OBUF2 REGF\[3\].RFW.BIT\[15\].FF/Q REGF\[3\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[15] sky130_fd_sc_hd__ebufn_2
Xfill_36_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[16\].RFW.BIT\[21\].OBUF2 REGF\[16\].RFW.BIT\[21\].FF/Q REGF\[16\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[21] sky130_fd_sc_hd__ebufn_2
Xfill_29_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[21\].RFW.BIT\[10\].OBUF2 REGF\[21\].RFW.BIT\[10\].FF/Q REGF\[21\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[10] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[5\].FF REGF\[27\].RFW.CG\[0\]/GCLK DW[5] VGND VGND VPWR VPWR
+ REGF\[27\].RFW.BIT\[5\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[26\].RFW.BIT\[7\].FF REGF\[26\].RFW.CG\[0\]/GCLK DW[7] VGND VGND VPWR VPWR
+ REGF\[26\].RFW.BIT\[7\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_23_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[17\].RFW.INV2\[2\] DEC1.D2.AND1/X VGND VGND VPWR VPWR REGF\[17\].RFW.INV2\[2\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_23_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_23_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_23_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.BIT\[24\].OBUF2 REGF\[12\].RFW.BIT\[24\].FF/Q REGF\[12\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[24] sky130_fd_sc_hd__ebufn_2
Xfill_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[25\].RFW.BIT\[9\].FF REGF\[25\].RFW.CG\[1\]/GCLK DW[9] VGND VGND VPWR VPWR
+ REGF\[25\].RFW.BIT\[9\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_48_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_48_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_48_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.BIT\[24\].FF REGF\[6\].RFW.CG\[3\]/GCLK DW[24] VGND VGND VPWR VPWR
+ REGF\[6\].RFW.BIT\[24\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[12\].RFW.BIT\[14\].FF REGF\[12\].RFW.CG\[1\]/GCLK DW[14] VGND VGND VPWR VPWR
+ REGF\[12\].RFW.BIT\[14\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_15_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgenblk1.RFW0.BIT\[25\].OBUF2 genblk1.RFW0.TIE\[7\]/LO genblk1.RFW0.INV2\[3\]/Y VGND
+ VGND VPWR VPWR DB[25] sky130_fd_sc_hd__ebufn_2
XDEC0.D2.ABUF\[1\] RA[1] VGND VGND VPWR VPWR DEC0.D2.AND7/B sky130_fd_sc_hd__clkbuf_2
XDEC0.D2.AND1 DEC0.D2.AND7/C DEC0.D2.AND7/B DEC0.D2.AND7/A DEC0.D2.AND7/D VGND VGND
+ VPWR VPWR DEC0.D2.AND1/X sky130_fd_sc_hd__and4bb_2
Xfill_41_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_34_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[20\].RFW.CGAND DEC2.D2.AND4/X WE VGND VGND VPWR VPWR REGF\[20\].RFW.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_27_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[23\].RFW.BIT\[24\].FF REGF\[23\].RFW.CG\[3\]/GCLK DW[24] VGND VGND VPWR VPWR
+ REGF\[23\].RFW.BIT\[24\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[13\].RFW.INV1\[3\] DEC0.D1.AND5/X VGND VGND VPWR VPWR REGF\[13\].RFW.INV1\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[11\].RFW.BIT\[12\].OBUF2 REGF\[11\].RFW.BIT\[12\].FF/Q REGF\[11\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[12] sky130_fd_sc_hd__ebufn_2
Xtap_56_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[9\].RFW.BIT\[8\].FF REGF\[9\].RFW.CG\[1\]/GCLK DW[8] VGND VGND VPWR VPWR REGF\[9\].RFW.BIT\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[9\].RFW.BIT\[27\].OBUF1 REGF\[9\].RFW.BIT\[27\].FF/Q REGF\[9\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[27] sky130_fd_sc_hd__ebufn_2
Xfill_18_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_18_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_18_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_62_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.BIT\[31\].FF REGF\[18\].RFW.CG\[3\]/GCLK DW[31] VGND VGND VPWR VPWR
+ REGF\[18\].RFW.BIT\[31\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[27\].RFW.BIT\[22\].OBUF1 REGF\[27\].RFW.BIT\[22\].FF/Q REGF\[27\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[22] sky130_fd_sc_hd__ebufn_2
Xfill_34_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_34_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_50_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_50_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_50_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_59_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_59_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_59_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_59_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_6_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_6_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_6_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_59_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_20_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_13_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[23\].RFW.BIT\[25\].OBUF1 REGF\[23\].RFW.BIT\[25\].FF/Q REGF\[23\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[25] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.INV2\[0\] DEC1.D0.AND4/X VGND VGND VPWR VPWR REGF\[4\].RFW.INV2\[0\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[8\].RFW.BIT\[15\].OBUF1 REGF\[8\].RFW.BIT\[15\].FF/Q REGF\[8\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[15] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[10\].OBUF1 REGF\[26\].RFW.BIT\[10\].FF/Q REGF\[26\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[10] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.BIT\[14\].FF REGF\[19\].RFW.CG\[1\]/GCLK DW[14] VGND VGND VPWR VPWR
+ REGF\[19\].RFW.BIT\[14\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[4\].RFW.CG\[2\] CLK REGF\[4\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[4\].RFW.CG\[2\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_54_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_20_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_20_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[27\].RFW.BIT\[26\].OBUF2 REGF\[27\].RFW.BIT\[26\].FF/Q REGF\[27\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[26] sky130_fd_sc_hd__ebufn_2
Xfill_20_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_29_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_29_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_29_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_29_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_29_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[4\].RFW.BIT\[18\].OBUF1 REGF\[4\].RFW.BIT\[18\].FF/Q REGF\[4\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[18] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[31\].OBUF1 REGF\[5\].RFW.BIT\[31\].FF/Q REGF\[5\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[31] sky130_fd_sc_hd__ebufn_2
Xfill_45_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_45_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[17\].RFW.BIT\[24\].OBUF1 REGF\[17\].RFW.BIT\[24\].FF/Q REGF\[17\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[24] sky130_fd_sc_hd__ebufn_2
Xfill_45_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_45_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_45_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_45_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_61_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_61_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_61_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_61_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[22\].RFW.BIT\[13\].OBUF1 REGF\[22\].RFW.BIT\[13\].FF/Q REGF\[22\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[13] sky130_fd_sc_hd__ebufn_2
Xfill_61_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_61_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDEC0.TIE VGND VGND VPWR VPWR DEC0.TIE/HI DEC0.TIE/LO sky130_fd_sc_hd__conb_1
XREGF\[10\].RFW.BIT\[0\].FF REGF\[10\].RFW.CG\[0\]/GCLK DW[0] VGND VGND VPWR VPWR
+ REGF\[10\].RFW.BIT\[0\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[23\].RFW.BIT\[29\].OBUF2 REGF\[23\].RFW.BIT\[29\].FF/Q REGF\[23\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[29] sky130_fd_sc_hd__ebufn_2
Xfill_9_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[8\].RFW.BIT\[19\].OBUF2 REGF\[8\].RFW.BIT\[19\].FF/Q REGF\[8\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[19] sky130_fd_sc_hd__ebufn_2
Xfill_11_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[4\].RFW.BIT\[15\].FF REGF\[4\].RFW.CG\[1\]/GCLK DW[15] VGND VGND VPWR VPWR
+ REGF\[4\].RFW.BIT\[15\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[13\].RFW.BIT\[27\].OBUF1 REGF\[13\].RFW.BIT\[27\].FF/Q REGF\[13\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[27] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[14\].OBUF2 REGF\[26\].RFW.BIT\[14\].FF/Q REGF\[26\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[14] sky130_fd_sc_hd__ebufn_2
Xtap_26_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[16\].RFW.BIT\[12\].OBUF1 REGF\[16\].RFW.BIT\[12\].FF/Q REGF\[16\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[12] sky130_fd_sc_hd__ebufn_2
Xfill_15_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_15_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_15_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_15_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_15_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[21\].RFW.BIT\[15\].FF REGF\[21\].RFW.CG\[1\]/GCLK DW[15] VGND VGND VPWR VPWR
+ REGF\[21\].RFW.BIT\[15\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_52_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_31_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_31_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_31_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.CG\[1\] CLK REGF\[18\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[18\].RFW.CG\[1\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_31_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[23\].RFW.BIT\[0\].FF REGF\[23\].RFW.CG\[0\]/GCLK DW[0] VGND VGND VPWR VPWR
+ REGF\[23\].RFW.BIT\[0\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_45_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[17\].RFW.BIT\[28\].OBUF2 REGF\[17\].RFW.BIT\[28\].FF/Q REGF\[17\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[28] sky130_fd_sc_hd__ebufn_2
Xtap_38_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[22\].RFW.BIT\[17\].OBUF2 REGF\[22\].RFW.BIT\[17\].FF/Q REGF\[22\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[17] sky130_fd_sc_hd__ebufn_2
XREGF\[23\].RFW.BIT\[30\].OBUF2 REGF\[23\].RFW.BIT\[30\].FF/Q REGF\[23\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[30] sky130_fd_sc_hd__ebufn_2
Xfill_56_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_56_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_56_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XREGF\[10\].RFW.BIT\[28\].FF REGF\[10\].RFW.CG\[3\]/GCLK DW[28] VGND VGND VPWR VPWR
+ REGF\[10\].RFW.BIT\[28\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[8\].RFW.BIT\[20\].OBUF2 REGF\[8\].RFW.BIT\[20\].FF/Q REGF\[8\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[20] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[22\].FF REGF\[16\].RFW.CG\[2\]/GCLK DW[22] VGND VGND VPWR VPWR
+ REGF\[16\].RFW.BIT\[22\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[22\].RFW.BIT\[2\].FF REGF\[22\].RFW.CG\[0\]/GCLK DW[2] VGND VGND VPWR VPWR
+ REGF\[22\].RFW.BIT\[2\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[12\].RFW.BIT\[15\].OBUF1 REGF\[12\].RFW.BIT\[15\].FF/Q REGF\[12\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[15] sky130_fd_sc_hd__ebufn_2
Xfill_59_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[15\].RFW.INV1\[0\] DEC0.D1.AND7/X VGND VGND VPWR VPWR REGF\[15\].RFW.INV1\[0\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[21\].RFW.BIT\[4\].FF REGF\[21\].RFW.CG\[0\]/GCLK DW[4] VGND VGND VPWR VPWR
+ REGF\[21\].RFW.BIT\[4\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_7_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XREGF\[30\].RFW.INV2\[1\] DEC1.D3.AND6/X VGND VGND VPWR VPWR REGF\[30\].RFW.INV2\[1\]/Y
+ sky130_fd_sc_hd__inv_4
Xgenblk1.RFW0.BIT\[16\].OBUF1 genblk1.RFW0.TIE\[2\]/LO genblk1.RFW0.INV1\[2\]/Y VGND
+ VGND VPWR VPWR DA[16] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.BIT\[23\].OBUF2 REGF\[4\].RFW.BIT\[23\].FF/Q REGF\[4\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[23] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[16\].OBUF2 REGF\[16\].RFW.BIT\[16\].FF/Q REGF\[16\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[16] sky130_fd_sc_hd__ebufn_2
XREGF\[20\].RFW.BIT\[6\].FF REGF\[20\].RFW.CG\[0\]/GCLK DW[6] VGND VGND VPWR VPWR
+ REGF\[20\].RFW.BIT\[6\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_24_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_26_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_26_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_26_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.BIT\[1\].FF REGF\[6\].RFW.CG\[0\]/GCLK DW[1] VGND VGND VPWR VPWR REGF\[6\].RFW.BIT\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[1\].RFW.BIT\[23\].FF REGF\[1\].RFW.CG\[2\]/GCLK DW[23] VGND VGND VPWR VPWR
+ REGF\[1\].RFW.BIT\[23\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_42_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_42_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_42_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[5\].RFW.BIT\[3\].FF REGF\[5\].RFW.CG\[0\]/GCLK DW[3] VGND VGND VPWR VPWR REGF\[5\].RFW.BIT\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[12\].RFW.BIT\[19\].OBUF2 REGF\[12\].RFW.BIT\[19\].FF/Q REGF\[12\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[19] sky130_fd_sc_hd__ebufn_2
Xfill_45_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_38_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[28\].RFW.BIT\[15\].FF REGF\[28\].RFW.CG\[1\]/GCLK DW[15] VGND VGND VPWR VPWR
+ REGF\[28\].RFW.BIT\[15\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[3\].RFW.BIT\[11\].OBUF2 REGF\[3\].RFW.BIT\[11\].FF/Q REGF\[3\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[11] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.BIT\[5\].FF REGF\[4\].RFW.CG\[0\]/GCLK DW[5] VGND VGND VPWR VPWR REGF\[4\].RFW.BIT\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[28\].RFW.BIT\[29\].OBUF1 REGF\[28\].RFW.BIT\[29\].FF/Q REGF\[28\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[29] sky130_fd_sc_hd__ebufn_2
Xfill_57_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[25\].RFW.INV2\[2\] DEC1.D3.AND1/X VGND VGND VPWR VPWR REGF\[25\].RFW.INV2\[2\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[17\].RFW.BIT\[28\].FF REGF\[17\].RFW.CG\[3\]/GCLK DW[28] VGND VGND VPWR VPWR
+ REGF\[17\].RFW.BIT\[28\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[13\].RFW.BIT\[30\].FF REGF\[13\].RFW.CG\[3\]/GCLK DW[30] VGND VGND VPWR VPWR
+ REGF\[13\].RFW.BIT\[30\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[3\].RFW.BIT\[7\].FF REGF\[3\].RFW.CG\[0\]/GCLK DW[7] VGND VGND VPWR VPWR REGF\[3\].RFW.BIT\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xfill_12_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_12_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_12_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_22_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.BIT\[20\].OBUF2 REGF\[12\].RFW.BIT\[20\].FF/Q REGF\[12\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[20] sky130_fd_sc_hd__ebufn_2
XREGF\[2\].RFW.BIT\[9\].FF REGF\[2\].RFW.CG\[1\]/GCLK DW[9] VGND VGND VPWR VPWR REGF\[2\].RFW.BIT\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xfill_37_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_37_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_37_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_37_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_37_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_53_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_53_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_53_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_53_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_53_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_53_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_9_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_9_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_9_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_9_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_9_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[27\].RFW.BIT\[17\].OBUF1 REGF\[27\].RFW.BIT\[17\].FF/Q REGF\[27\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[17] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.BIT\[30\].OBUF1 REGF\[28\].RFW.BIT\[30\].FF/Q REGF\[28\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[30] sky130_fd_sc_hd__ebufn_2
Xfill_50_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[21\].RFW.INV1\[3\] DEC0.D2.AND5/X VGND VGND VPWR VPWR REGF\[21\].RFW.INV1\[3\]/Y
+ sky130_fd_sc_hd__inv_4
Xgenblk1.RFW0.BIT\[21\].OBUF2 genblk1.RFW0.TIE\[6\]/LO genblk1.RFW0.INV2\[2\]/Y VGND
+ VGND VPWR VPWR DB[21] sky130_fd_sc_hd__ebufn_2
Xfill_43_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_36_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_29_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[2\].RFW.BIT\[29\].FF REGF\[2\].RFW.CG\[3\]/GCLK DW[29] VGND VGND VPWR VPWR
+ REGF\[2\].RFW.BIT\[29\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[8\].RFW.BIT\[23\].FF REGF\[8\].RFW.CG\[2\]/GCLK DW[23] VGND VGND VPWR VPWR
+ REGF\[8\].RFW.BIT\[23\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[14\].RFW.BIT\[13\].FF REGF\[14\].RFW.CG\[1\]/GCLK DW[13] VGND VGND VPWR VPWR
+ REGF\[14\].RFW.BIT\[13\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[30\].RFW.BIT\[16\].FF REGF\[30\].RFW.CG\[2\]/GCLK DW[16] VGND VGND VPWR VPWR
+ REGF\[30\].RFW.BIT\[16\].FF/Q sky130_fd_sc_hd__dfxtp_1
XDEC1.D1.AND0 DEC1.D1.AND7/A DEC1.D1.AND7/B DEC1.D1.AND7/C DEC1.D1.AND7/D VGND VGND
+ VPWR VPWR DEC1.D1.AND0/Y sky130_fd_sc_hd__nor4b_2
XREGF\[9\].RFW.BIT\[23\].OBUF1 REGF\[9\].RFW.BIT\[23\].FF/Q REGF\[9\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[23] sky130_fd_sc_hd__ebufn_2
Xfill_23_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_23_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_23_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_23_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_23_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[25\].RFW.BIT\[23\].FF REGF\[25\].RFW.CG\[2\]/GCLK DW[23] VGND VGND VPWR VPWR
+ REGF\[25\].RFW.BIT\[23\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[11\].RFW.BIT\[9\].OBUF1 REGF\[11\].RFW.BIT\[9\].FF/Q REGF\[11\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[9] sky130_fd_sc_hd__ebufn_2
Xtap_20_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_48_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_48_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_48_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[1\].RFW.BIT\[8\].OBUF1 REGF\[1\].RFW.BIT\[8\].FF/Q REGF\[1\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[8] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[26\].OBUF1 REGF\[5\].RFW.BIT\[26\].FF/Q REGF\[5\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[26] sky130_fd_sc_hd__ebufn_2
XDEC0.D2.AND2 DEC0.D2.AND7/C DEC0.D2.AND7/A DEC0.D2.AND7/B DEC0.D2.AND7/D VGND VGND
+ VPWR VPWR DEC0.D2.AND2/X sky130_fd_sc_hd__and4bb_2
XREGF\[27\].RFW.CG\[3\] CLK REGF\[27\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[27\].RFW.CG\[3\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[17\].RFW.BIT\[19\].OBUF1 REGF\[17\].RFW.BIT\[19\].FF/Q REGF\[17\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[19] sky130_fd_sc_hd__ebufn_2
XREGF\[23\].RFW.BIT\[21\].OBUF1 REGF\[23\].RFW.BIT\[21\].FF/Q REGF\[23\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[21] sky130_fd_sc_hd__ebufn_2
Xfill_41_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_27_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[8\].RFW.BIT\[11\].OBUF1 REGF\[8\].RFW.BIT\[11\].FF/Q REGF\[8\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[11] sky130_fd_sc_hd__ebufn_2
Xfill_1_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[13\].RFW.BIT\[9\].OBUF1 REGF\[13\].RFW.BIT\[9\].FF/Q REGF\[13\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[9] sky130_fd_sc_hd__ebufn_2
Xtap_56_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[9\].RFW.BIT\[27\].OBUF2 REGF\[9\].RFW.BIT\[27\].FF/Q REGF\[9\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[27] sky130_fd_sc_hd__ebufn_2
XDEC0.D0.ABUF\[0\] RA[0] VGND VGND VPWR VPWR DEC0.D0.AND7/A sky130_fd_sc_hd__clkbuf_2
XREGF\[26\].RFW.CG\[0\] CLK REGF\[26\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[26\].RFW.CG\[0\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[1\].RFW.BIT\[29\].OBUF1 REGF\[1\].RFW.BIT\[29\].FF/Q REGF\[1\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[29] sky130_fd_sc_hd__ebufn_2
Xfill_18_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_18_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_18_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[3\].RFW.BIT\[8\].OBUF1 REGF\[3\].RFW.BIT\[8\].FF/Q REGF\[3\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[8] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[22\].OBUF2 REGF\[27\].RFW.BIT\[22\].FF/Q REGF\[27\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[22] sky130_fd_sc_hd__ebufn_2
Xfill_34_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_34_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_34_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[9\].RFW.BIT\[29\].FF REGF\[9\].RFW.CG\[3\]/GCLK DW[29] VGND VGND VPWR VPWR
+ REGF\[9\].RFW.BIT\[29\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[15\].RFW.BIT\[19\].FF REGF\[15\].RFW.CG\[2\]/GCLK DW[19] VGND VGND VPWR VPWR
+ REGF\[15\].RFW.BIT\[19\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[5\].RFW.BIT\[31\].FF REGF\[5\].RFW.CG\[3\]/GCLK DW[31] VGND VGND VPWR VPWR
+ REGF\[5\].RFW.BIT\[31\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[11\].RFW.BIT\[21\].FF REGF\[11\].RFW.CG\[2\]/GCLK DW[21] VGND VGND VPWR VPWR
+ REGF\[11\].RFW.BIT\[21\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_50_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_50_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_50_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[4\].RFW.BIT\[14\].OBUF1 REGF\[4\].RFW.BIT\[14\].FF/Q REGF\[4\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[14] sky130_fd_sc_hd__ebufn_2
Xfill_59_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[17\].RFW.BIT\[20\].OBUF1 REGF\[17\].RFW.BIT\[20\].FF/Q REGF\[17\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[20] sky130_fd_sc_hd__ebufn_2
Xfill_59_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_59_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_59_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_59_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_6_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_6_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_6_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_59_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[7\].RFW.INV2\[1\] DEC1.D0.AND7/X VGND VGND VPWR VPWR REGF\[7\].RFW.INV2\[1\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[15\].RFW.BIT\[9\].OBUF1 REGF\[15\].RFW.BIT\[9\].FF/Q REGF\[15\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[9] sky130_fd_sc_hd__ebufn_2
Xfill_20_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_13_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[15\].RFW.CG\[3\] CLK REGF\[15\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[15\].RFW.CG\[3\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[23\].RFW.BIT\[25\].OBUF2 REGF\[23\].RFW.BIT\[25\].FF/Q REGF\[23\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[25] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[29\].FF REGF\[26\].RFW.CG\[3\]/GCLK DW[29] VGND VGND VPWR VPWR
+ REGF\[26\].RFW.BIT\[29\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[22\].RFW.BIT\[31\].FF REGF\[22\].RFW.CG\[3\]/GCLK DW[31] VGND VGND VPWR VPWR
+ REGF\[22\].RFW.BIT\[31\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[8\].RFW.BIT\[15\].OBUF2 REGF\[8\].RFW.BIT\[15\].FF/Q REGF\[8\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[15] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[8\].OBUF1 REGF\[5\].RFW.BIT\[8\].FF/Q REGF\[5\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[8] sky130_fd_sc_hd__ebufn_2
XREGF\[1\].RFW.BIT\[30\].OBUF1 REGF\[1\].RFW.BIT\[30\].FF/Q REGF\[1\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[30] sky130_fd_sc_hd__ebufn_2
XREGF\[13\].RFW.BIT\[23\].OBUF1 REGF\[13\].RFW.BIT\[23\].FF/Q REGF\[13\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[23] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[10\].OBUF2 REGF\[26\].RFW.BIT\[10\].FF/Q REGF\[26\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[10] sky130_fd_sc_hd__ebufn_2
XREGF\[14\].RFW.CG\[0\] CLK REGF\[14\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[14\].RFW.CG\[0\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_54_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.BIT\[14\].FF REGF\[6\].RFW.CG\[1\]/GCLK DW[14] VGND VGND VPWR VPWR
+ REGF\[6\].RFW.BIT\[14\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_20_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_20_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XREGF\[3\].RFW.INV1\[2\] DEC0.D0.AND3/X VGND VGND VPWR VPWR REGF\[3\].RFW.INV1\[2\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[17\].RFW.BIT\[9\].OBUF1 REGF\[17\].RFW.BIT\[9\].FF/Q REGF\[17\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[9] sky130_fd_sc_hd__ebufn_2
Xfill_29_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_29_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_29_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_29_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[4\].RFW.BIT\[18\].OBUF2 REGF\[4\].RFW.BIT\[18\].FF/Q REGF\[4\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[18] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[31\].OBUF2 REGF\[5\].RFW.BIT\[31\].FF/Q REGF\[5\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[31] sky130_fd_sc_hd__ebufn_2
Xfill_45_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_45_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_45_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_45_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_45_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[17\].RFW.BIT\[24\].OBUF2 REGF\[17\].RFW.BIT\[24\].FF/Q REGF\[17\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[24] sky130_fd_sc_hd__ebufn_2
Xfill_61_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_61_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_61_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_61_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XREGF\[7\].RFW.BIT\[8\].OBUF1 REGF\[7\].RFW.BIT\[8\].FF/Q REGF\[7\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[8] sky130_fd_sc_hd__ebufn_2
XREGF\[22\].RFW.BIT\[13\].OBUF2 REGF\[22\].RFW.BIT\[13\].FF/Q REGF\[22\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[13] sky130_fd_sc_hd__ebufn_2
Xfill_61_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_61_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[23\].RFW.INV1\[0\] DEC0.D2.AND7/X VGND VGND VPWR VPWR REGF\[23\].RFW.INV1\[0\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[10\].RFW.BIT\[7\].OBUF1 REGF\[10\].RFW.BIT\[7\].FF/Q REGF\[10\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[7] sky130_fd_sc_hd__ebufn_2
XREGF\[23\].RFW.BIT\[14\].FF REGF\[23\].RFW.CG\[1\]/GCLK DW[14] VGND VGND VPWR VPWR
+ REGF\[23\].RFW.BIT\[14\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[12\].RFW.BIT\[11\].OBUF1 REGF\[12\].RFW.BIT\[11\].FF/Q REGF\[12\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[11] sky130_fd_sc_hd__ebufn_2
Xfill_9_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_11_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.BIT\[27\].FF REGF\[12\].RFW.CG\[3\]/GCLK DW[27] VGND VGND VPWR VPWR
+ REGF\[12\].RFW.BIT\[27\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[19\].RFW.BIT\[9\].OBUF1 REGF\[19\].RFW.BIT\[9\].FF/Q REGF\[19\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[9] sky130_fd_sc_hd__ebufn_2
XREGF\[13\].RFW.BIT\[27\].OBUF2 REGF\[13\].RFW.BIT\[27\].FF/Q REGF\[13\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[27] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.BIT\[21\].FF REGF\[18\].RFW.CG\[2\]/GCLK DW[21] VGND VGND VPWR VPWR
+ REGF\[18\].RFW.BIT\[21\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[9\].RFW.BIT\[8\].OBUF1 REGF\[9\].RFW.BIT\[8\].FF/Q REGF\[9\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[8] sky130_fd_sc_hd__ebufn_2
Xgenblk1.RFW0.BIT\[12\].OBUF1 genblk1.RFW0.TIE\[1\]/LO genblk1.RFW0.INV1\[1\]/Y VGND
+ VGND VPWR VPWR DA[12] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[12\].OBUF2 REGF\[16\].RFW.BIT\[12\].FF/Q REGF\[16\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[12] sky130_fd_sc_hd__ebufn_2
Xfill_15_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_15_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_15_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_15_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.BIT\[7\].OBUF1 REGF\[12\].RFW.BIT\[7\].FF/Q REGF\[12\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[7] sky130_fd_sc_hd__ebufn_2
Xfill_15_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_31_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_31_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_31_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_52_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_31_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_31_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_45_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_38_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[29\].RFW.BIT\[31\].FF REGF\[29\].RFW.CG\[3\]/GCLK DW[31] VGND VGND VPWR VPWR
+ REGF\[29\].RFW.BIT\[31\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[2\].RFW.BIT\[6\].OBUF1 REGF\[2\].RFW.BIT\[6\].FF/Q REGF\[2\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[6] sky130_fd_sc_hd__ebufn_2
Xfill_56_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_56_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_56_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[18\].RFW.INV1\[1\] DEC0.D2.AND2/X VGND VGND VPWR VPWR REGF\[18\].RFW.INV1\[1\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[12\].RFW.BIT\[15\].OBUF2 REGF\[12\].RFW.BIT\[15\].FF/Q REGF\[12\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[15] sky130_fd_sc_hd__ebufn_2
XREGF\[3\].RFW.BIT\[22\].FF REGF\[3\].RFW.CG\[2\]/GCLK DW[22] VGND VGND VPWR VPWR
+ REGF\[3\].RFW.BIT\[22\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[30\].RFW.BIT\[29\].OBUF1 REGF\[30\].RFW.BIT\[29\].FF/Q REGF\[30\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[29] sky130_fd_sc_hd__ebufn_2
Xgenblk1.RFW0.TIE\[2\] VGND VGND VPWR VPWR genblk1.RFW0.TIE\[2\]/HI genblk1.RFW0.TIE\[2\]/LO
+ sky130_fd_sc_hd__conb_1
Xfill_59_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[14\].RFW.BIT\[7\].OBUF1 REGF\[14\].RFW.BIT\[7\].FF/Q REGF\[14\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[7] sky130_fd_sc_hd__ebufn_2
Xfill_7_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[28\].RFW.BIT\[25\].OBUF1 REGF\[28\].RFW.BIT\[25\].FF/Q REGF\[28\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[25] sky130_fd_sc_hd__ebufn_2
Xgenblk1.RFW0.BIT\[16\].OBUF2 genblk1.RFW0.TIE\[6\]/LO genblk1.RFW0.INV2\[2\]/Y VGND
+ VGND VPWR VPWR DB[16] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.BIT\[6\].OBUF1 REGF\[4\].RFW.BIT\[6\].FF/Q REGF\[4\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[6] sky130_fd_sc_hd__ebufn_2
XREGF\[20\].RFW.BIT\[22\].FF REGF\[20\].RFW.CG\[2\]/GCLK DW[22] VGND VGND VPWR VPWR
+ REGF\[20\].RFW.BIT\[22\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_24_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_26_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_26_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_26_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_42_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_42_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_42_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[24\].RFW.BIT\[28\].OBUF1 REGF\[24\].RFW.BIT\[28\].FF/Q REGF\[24\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[28] sky130_fd_sc_hd__ebufn_2
Xtap_50_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[19\].RFW.BIT\[27\].FF REGF\[19\].RFW.CG\[3\]/GCLK DW[27] VGND VGND VPWR VPWR
+ REGF\[19\].RFW.BIT\[27\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[16\].RFW.BIT\[7\].OBUF1 REGF\[16\].RFW.BIT\[7\].FF/Q REGF\[16\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[7] sky130_fd_sc_hd__ebufn_2
XREGF\[30\].RFW.BIT\[30\].OBUF1 REGF\[30\].RFW.BIT\[30\].FF/Q REGF\[30\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[30] sky130_fd_sc_hd__ebufn_2
XREGF\[9\].RFW.BIT\[18\].OBUF1 REGF\[9\].RFW.BIT\[18\].FF/Q REGF\[9\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[18] sky130_fd_sc_hd__ebufn_2
Xfill_38_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[27\].RFW.BIT\[13\].OBUF1 REGF\[27\].RFW.BIT\[13\].FF/Q REGF\[27\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[13] sky130_fd_sc_hd__ebufn_2
XREGF\[6\].RFW.BIT\[6\].OBUF1 REGF\[6\].RFW.BIT\[6\].FF/Q REGF\[6\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[6] sky130_fd_sc_hd__ebufn_2
XREGF\[12\].RFW.INV2\[2\] DEC1.D1.AND4/X VGND VGND VPWR VPWR REGF\[12\].RFW.INV2\[2\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[28\].RFW.INV2\[3\] DEC1.D3.AND4/X VGND VGND VPWR VPWR REGF\[28\].RFW.INV2\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[28\].RFW.BIT\[29\].OBUF2 REGF\[28\].RFW.BIT\[29\].FF/Q REGF\[28\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[29] sky130_fd_sc_hd__ebufn_2
Xfill_57_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_5_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.BIT\[27\].OBUF1 REGF\[18\].RFW.BIT\[27\].FF/Q REGF\[18\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[27] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.BIT\[7\].OBUF1 REGF\[18\].RFW.BIT\[7\].FF/Q REGF\[18\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[7] sky130_fd_sc_hd__ebufn_2
XREGF\[23\].RFW.BIT\[16\].OBUF1 REGF\[23\].RFW.BIT\[16\].FF/Q REGF\[23\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[16] sky130_fd_sc_hd__ebufn_2
Xfill_12_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_12_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[10\].RFW.BIT\[18\].FF REGF\[10\].RFW.CG\[2\]/GCLK DW[18] VGND VGND VPWR VPWR
+ REGF\[10\].RFW.BIT\[18\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_12_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XREGF\[4\].RFW.BIT\[28\].FF REGF\[4\].RFW.CG\[3\]/GCLK DW[28] VGND VGND VPWR VPWR
+ REGF\[4\].RFW.BIT\[28\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[16\].RFW.BIT\[12\].FF REGF\[16\].RFW.CG\[1\]/GCLK DW[12] VGND VGND VPWR VPWR
+ REGF\[16\].RFW.BIT\[12\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_22_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_15_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[8\].RFW.BIT\[6\].OBUF1 REGF\[8\].RFW.BIT\[6\].FF/Q REGF\[8\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[6] sky130_fd_sc_hd__ebufn_2
Xfill_37_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_37_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_37_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_37_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_37_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_53_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_53_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_53_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_53_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[11\].RFW.BIT\[5\].OBUF1 REGF\[11\].RFW.BIT\[5\].FF/Q REGF\[11\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[5] sky130_fd_sc_hd__ebufn_2
Xfill_53_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_9_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[23\].RFW.CG\[2\] CLK REGF\[23\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[23\].RFW.CG\[2\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_9_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_9_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_9_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[21\].RFW.BIT\[28\].FF REGF\[21\].RFW.CG\[3\]/GCLK DW[28] VGND VGND VPWR VPWR
+ REGF\[21\].RFW.BIT\[28\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[27\].RFW.BIT\[17\].OBUF2 REGF\[27\].RFW.BIT\[17\].FF/Q REGF\[27\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[17] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.BIT\[30\].OBUF2 REGF\[28\].RFW.BIT\[30\].FF/Q REGF\[28\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[30] sky130_fd_sc_hd__ebufn_2
XREGF\[1\].RFW.BIT\[4\].OBUF1 REGF\[1\].RFW.BIT\[4\].FF/Q REGF\[1\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[4] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[22\].FF REGF\[27\].RFW.CG\[2\]/GCLK DW[22] VGND VGND VPWR VPWR
+ REGF\[27\].RFW.BIT\[22\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_50_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_43_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_36_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[5\].RFW.BIT\[22\].OBUF1 REGF\[5\].RFW.BIT\[22\].FF/Q REGF\[5\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[22] sky130_fd_sc_hd__ebufn_2
Xfill_29_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[17\].RFW.BIT\[15\].OBUF1 REGF\[17\].RFW.BIT\[15\].FF/Q REGF\[17\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[15] sky130_fd_sc_hd__ebufn_2
XREGF\[1\].RFW.BIT\[13\].FF REGF\[1\].RFW.CG\[1\]/GCLK DW[13] VGND VGND VPWR VPWR
+ REGF\[1\].RFW.BIT\[13\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[13\].RFW.BIT\[5\].OBUF1 REGF\[13\].RFW.BIT\[5\].FF/Q REGF\[13\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[5] sky130_fd_sc_hd__ebufn_2
XDEC1.D1.AND1 DEC1.D1.AND7/C DEC1.D1.AND7/B DEC1.D1.AND7/A DEC1.D1.AND7/D VGND VGND
+ VPWR VPWR DEC1.D1.AND1/X sky130_fd_sc_hd__and4bb_2
XREGF\[9\].RFW.BIT\[23\].OBUF2 REGF\[9\].RFW.BIT\[23\].FF/Q REGF\[9\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[23] sky130_fd_sc_hd__ebufn_2
Xfill_23_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_23_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_23_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[1\].RFW.BIT\[25\].OBUF1 REGF\[1\].RFW.BIT\[25\].FF/Q REGF\[1\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[25] sky130_fd_sc_hd__ebufn_2
Xfill_23_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_23_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.BIT\[4\].OBUF1 REGF\[3\].RFW.BIT\[4\].FF/Q REGF\[3\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[4] sky130_fd_sc_hd__ebufn_2
XREGF\[14\].RFW.BIT\[31\].OBUF1 REGF\[14\].RFW.BIT\[31\].FF/Q REGF\[14\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[31] sky130_fd_sc_hd__ebufn_2
XREGF\[13\].RFW.BIT\[18\].OBUF1 REGF\[13\].RFW.BIT\[18\].FF/Q REGF\[13\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[18] sky130_fd_sc_hd__ebufn_2
XREGF\[11\].RFW.BIT\[9\].OBUF2 REGF\[11\].RFW.BIT\[9\].FF/Q REGF\[11\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[9] sky130_fd_sc_hd__ebufn_2
Xtap_20_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_48_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_48_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_48_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[4\].RFW.BIT\[10\].OBUF1 REGF\[4\].RFW.BIT\[10\].FF/Q REGF\[4\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[10] sky130_fd_sc_hd__ebufn_2
XREGF\[11\].RFW.CG\[2\] CLK REGF\[11\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[11\].RFW.CG\[2\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[1\].RFW.BIT\[8\].OBUF2 REGF\[1\].RFW.BIT\[8\].FF/Q REGF\[1\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[8] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[26\].OBUF2 REGF\[5\].RFW.BIT\[26\].FF/Q REGF\[5\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[26] sky130_fd_sc_hd__ebufn_2
XDEC0.D2.AND3 DEC0.D2.AND7/C DEC0.D2.AND7/B DEC0.D2.AND7/A DEC0.D2.AND7/D VGND VGND
+ VPWR VPWR DEC0.D2.AND3/X sky130_fd_sc_hd__and4b_2
XREGF\[15\].RFW.BIT\[5\].OBUF1 REGF\[15\].RFW.BIT\[5\].FF/Q REGF\[15\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[5] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.BIT\[18\].FF REGF\[17\].RFW.CG\[2\]/GCLK DW[18] VGND VGND VPWR VPWR
+ REGF\[17\].RFW.BIT\[18\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[17\].RFW.BIT\[19\].OBUF2 REGF\[17\].RFW.BIT\[19\].FF/Q REGF\[17\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[19] sky130_fd_sc_hd__ebufn_2
XREGF\[7\].RFW.BIT\[30\].FF REGF\[7\].RFW.CG\[3\]/GCLK DW[30] VGND VGND VPWR VPWR
+ REGF\[7\].RFW.BIT\[30\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[13\].RFW.BIT\[20\].FF REGF\[13\].RFW.CG\[2\]/GCLK DW[20] VGND VGND VPWR VPWR
+ REGF\[13\].RFW.BIT\[20\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[23\].RFW.BIT\[21\].OBUF2 REGF\[23\].RFW.BIT\[21\].FF/Q REGF\[23\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[21] sky130_fd_sc_hd__ebufn_2
Xfill_41_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[5\].RFW.BIT\[4\].OBUF1 REGF\[5\].RFW.BIT\[4\].FF/Q REGF\[5\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[4] sky130_fd_sc_hd__ebufn_2
Xfill_27_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XREGF\[8\].RFW.BIT\[11\].OBUF2 REGF\[8\].RFW.BIT\[11\].FF/Q REGF\[8\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[11] sky130_fd_sc_hd__ebufn_2
Xfill_1_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[13\].RFW.BIT\[9\].OBUF2 REGF\[13\].RFW.BIT\[9\].FF/Q REGF\[13\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[9] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.BIT\[28\].FF REGF\[28\].RFW.CG\[3\]/GCLK DW[28] VGND VGND VPWR VPWR
+ REGF\[28\].RFW.BIT\[28\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[1\].RFW.BIT\[29\].OBUF2 REGF\[1\].RFW.BIT\[29\].FF/Q REGF\[1\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[29] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[30\].FF REGF\[24\].RFW.CG\[3\]/GCLK DW[30] VGND VGND VPWR VPWR
+ REGF\[24\].RFW.BIT\[30\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_18_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_18_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.BIT\[8\].OBUF2 REGF\[3\].RFW.BIT\[8\].FF/Q REGF\[3\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[8] sky130_fd_sc_hd__ebufn_2
Xfill_18_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_34_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[17\].RFW.BIT\[5\].OBUF1 REGF\[17\].RFW.BIT\[5\].FF/Q REGF\[17\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[5] sky130_fd_sc_hd__ebufn_2
Xfill_34_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.INV1\[0\] DEC0.D3.AND7/X VGND VGND VPWR VPWR REGF\[31\].RFW.INV1\[0\]/Y
+ sky130_fd_sc_hd__inv_4
Xgenblk1.RFW0.BIT\[9\].OBUF1 genblk1.RFW0.TIE\[1\]/LO genblk1.RFW0.INV1\[1\]/Y VGND
+ VGND VPWR VPWR DA[9] sky130_fd_sc_hd__ebufn_2
Xfill_50_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_50_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[4\].RFW.BIT\[14\].OBUF2 REGF\[4\].RFW.BIT\[14\].FF/Q REGF\[4\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[14] sky130_fd_sc_hd__ebufn_2
Xfill_50_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_59_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XREGF\[17\].RFW.BIT\[20\].OBUF2 REGF\[17\].RFW.BIT\[20\].FF/Q REGF\[17\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[20] sky130_fd_sc_hd__ebufn_2
Xfill_59_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_59_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_59_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_6_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_6_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[2\].RFW.BIT\[19\].FF REGF\[2\].RFW.CG\[2\]/GCLK DW[19] VGND VGND VPWR VPWR
+ REGF\[2\].RFW.BIT\[19\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_59_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_59_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[7\].RFW.BIT\[4\].OBUF1 REGF\[7\].RFW.BIT\[4\].FF/Q REGF\[7\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[4] sky130_fd_sc_hd__ebufn_2
XREGF\[8\].RFW.BIT\[13\].FF REGF\[8\].RFW.CG\[1\]/GCLK DW[13] VGND VGND VPWR VPWR
+ REGF\[8\].RFW.BIT\[13\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[15\].RFW.BIT\[9\].OBUF2 REGF\[15\].RFW.BIT\[9\].FF/Q REGF\[15\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[9] sky130_fd_sc_hd__ebufn_2
Xfill_20_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[10\].RFW.BIT\[3\].OBUF1 REGF\[10\].RFW.BIT\[3\].FF/Q REGF\[10\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[3] sky130_fd_sc_hd__ebufn_2
Xfill_13_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[5\].RFW.BIT\[8\].OBUF2 REGF\[5\].RFW.BIT\[8\].FF/Q REGF\[5\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[8] sky130_fd_sc_hd__ebufn_2
XREGF\[1\].RFW.BIT\[30\].OBUF2 REGF\[1\].RFW.BIT\[30\].FF/Q REGF\[1\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[30] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.BIT\[5\].OBUF1 REGF\[19\].RFW.BIT\[5\].FF/Q REGF\[19\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[5] sky130_fd_sc_hd__ebufn_2
XREGF\[13\].RFW.BIT\[23\].OBUF2 REGF\[13\].RFW.BIT\[23\].FF/Q REGF\[13\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[23] sky130_fd_sc_hd__ebufn_2
Xfill_32_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[25\].RFW.BIT\[13\].FF REGF\[25\].RFW.CG\[1\]/GCLK DW[13] VGND VGND VPWR VPWR
+ REGF\[25\].RFW.BIT\[13\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[6\].RFW.INV1\[3\] DEC0.D0.AND6/X VGND VGND VPWR VPWR REGF\[6\].RFW.INV1\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[9\].RFW.BIT\[4\].OBUF1 REGF\[9\].RFW.BIT\[4\].FF/Q REGF\[9\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[4] sky130_fd_sc_hd__ebufn_2
Xtap_54_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_20_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.BIT\[0\].FF REGF\[18\].RFW.CG\[0\]/GCLK DW[0] VGND VGND VPWR VPWR
+ REGF\[18\].RFW.BIT\[0\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_20_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[10\].RFW.INV1\[0\] DEC0.D1.AND2/X VGND VGND VPWR VPWR REGF\[10\].RFW.INV1\[0\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[14\].RFW.BIT\[26\].FF REGF\[14\].RFW.CG\[3\]/GCLK DW[26] VGND VGND VPWR VPWR
+ REGF\[14\].RFW.BIT\[26\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[17\].RFW.BIT\[9\].OBUF2 REGF\[17\].RFW.BIT\[9\].FF/Q REGF\[17\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[9] sky130_fd_sc_hd__ebufn_2
XREGF\[12\].RFW.BIT\[3\].OBUF1 REGF\[12\].RFW.BIT\[3\].FF/Q REGF\[12\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[3] sky130_fd_sc_hd__ebufn_2
Xfill_29_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_29_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_29_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[30\].RFW.BIT\[29\].FF REGF\[30\].RFW.CG\[3\]/GCLK DW[29] VGND VGND VPWR VPWR
+ REGF\[30\].RFW.BIT\[29\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_29_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_29_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[26\].RFW.INV1\[1\] DEC0.D3.AND2/X VGND VGND VPWR VPWR REGF\[26\].RFW.INV1\[1\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_45_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_45_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_45_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_45_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_45_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_61_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_61_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_61_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[7\].RFW.BIT\[8\].OBUF2 REGF\[7\].RFW.BIT\[8\].FF/Q REGF\[7\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[8] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.BIT\[2\].FF REGF\[17\].RFW.CG\[0\]/GCLK DW[2] VGND VGND VPWR VPWR
+ REGF\[17\].RFW.BIT\[2\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[2\].RFW.BIT\[2\].OBUF1 REGF\[2\].RFW.BIT\[2\].FF/Q REGF\[2\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[2] sky130_fd_sc_hd__ebufn_2
Xfill_61_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_61_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[10\].RFW.BIT\[7\].OBUF2 REGF\[10\].RFW.BIT\[7\].FF/Q REGF\[10\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[7] sky130_fd_sc_hd__ebufn_2
XREGF\[12\].RFW.BIT\[11\].OBUF2 REGF\[12\].RFW.BIT\[11\].FF/Q REGF\[12\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[11] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[4\].FF REGF\[16\].RFW.CG\[0\]/GCLK DW[4] VGND VGND VPWR VPWR
+ REGF\[16\].RFW.BIT\[4\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_11_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_9_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[30\].RFW.BIT\[25\].OBUF1 REGF\[30\].RFW.BIT\[25\].FF/Q REGF\[30\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[25] sky130_fd_sc_hd__ebufn_2
XREGF\[14\].RFW.BIT\[3\].OBUF1 REGF\[14\].RFW.BIT\[3\].FF/Q REGF\[14\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[3] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.BIT\[9\].OBUF2 REGF\[19\].RFW.BIT\[9\].FF/Q REGF\[19\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[9] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.BIT\[21\].OBUF1 REGF\[28\].RFW.BIT\[21\].FF/Q REGF\[28\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[21] sky130_fd_sc_hd__ebufn_2
XREGF\[15\].RFW.BIT\[6\].FF REGF\[15\].RFW.CG\[0\]/GCLK DW[6] VGND VGND VPWR VPWR
+ REGF\[15\].RFW.BIT\[6\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_7_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[9\].RFW.BIT\[19\].FF REGF\[9\].RFW.CG\[2\]/GCLK DW[19] VGND VGND VPWR VPWR
+ REGF\[9\].RFW.BIT\[19\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[9\].RFW.BIT\[8\].OBUF2 REGF\[9\].RFW.BIT\[8\].FF/Q REGF\[9\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[8] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[21\].FF REGF\[5\].RFW.CG\[2\]/GCLK DW[21] VGND VGND VPWR VPWR
+ REGF\[5\].RFW.BIT\[21\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[11\].RFW.BIT\[11\].FF REGF\[11\].RFW.CG\[1\]/GCLK DW[11] VGND VGND VPWR VPWR
+ REGF\[11\].RFW.BIT\[11\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xgenblk1.RFW0.BIT\[12\].OBUF2 genblk1.RFW0.TIE\[5\]/LO genblk1.RFW0.INV2\[1\]/Y VGND
+ VGND VPWR VPWR DB[12] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.BIT\[2\].OBUF1 REGF\[4\].RFW.BIT\[2\].FF/Q REGF\[4\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[2] sky130_fd_sc_hd__ebufn_2
Xfill_15_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_15_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_15_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.BIT\[7\].OBUF2 REGF\[12\].RFW.BIT\[7\].FF/Q REGF\[12\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[7] sky130_fd_sc_hd__ebufn_2
XREGF\[14\].RFW.BIT\[8\].FF REGF\[14\].RFW.CG\[1\]/GCLK DW[8] VGND VGND VPWR VPWR
+ REGF\[14\].RFW.BIT\[8\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_31_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_31_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xtap_52_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_31_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_31_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_31_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_45_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.BIT\[29\].OBUF1 REGF\[6\].RFW.BIT\[29\].FF/Q REGF\[6\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[29] sky130_fd_sc_hd__ebufn_2
Xtap_38_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.CG\[1\] CLK REGF\[31\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[31\].RFW.CG\[1\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[2\].RFW.BIT\[6\].OBUF2 REGF\[2\].RFW.BIT\[6\].FF/Q REGF\[2\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[6] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.BIT\[4\].FF REGF\[29\].RFW.CG\[0\]/GCLK DW[4] VGND VGND VPWR VPWR
+ REGF\[29\].RFW.BIT\[4\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_56_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_56_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[24\].RFW.BIT\[24\].OBUF1 REGF\[24\].RFW.BIT\[24\].FF/Q REGF\[24\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[24] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[19\].FF REGF\[26\].RFW.CG\[2\]/GCLK DW[19] VGND VGND VPWR VPWR
+ REGF\[26\].RFW.BIT\[19\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_56_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.INV2\[2\] DEC1.D2.AND4/X VGND VGND VPWR VPWR REGF\[20\].RFW.INV2\[2\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[22\].RFW.BIT\[21\].FF REGF\[22\].RFW.CG\[2\]/GCLK DW[21] VGND VGND VPWR VPWR
+ REGF\[22\].RFW.BIT\[21\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[16\].RFW.BIT\[3\].OBUF1 REGF\[16\].RFW.BIT\[3\].FF/Q REGF\[16\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[3] sky130_fd_sc_hd__ebufn_2
XREGF\[9\].RFW.BIT\[14\].OBUF1 REGF\[9\].RFW.BIT\[14\].FF/Q REGF\[9\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[14] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.BIT\[6\].FF REGF\[28\].RFW.CG\[0\]/GCLK DW[6] VGND VGND VPWR VPWR
+ REGF\[28\].RFW.BIT\[6\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[6\].RFW.BIT\[2\].OBUF1 REGF\[6\].RFW.BIT\[2\].FF/Q REGF\[6\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[2] sky130_fd_sc_hd__ebufn_2
XREGF\[30\].RFW.BIT\[29\].OBUF2 REGF\[30\].RFW.BIT\[29\].FF/Q REGF\[30\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[29] sky130_fd_sc_hd__ebufn_2
Xfill_59_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[14\].RFW.BIT\[7\].OBUF2 REGF\[14\].RFW.BIT\[7\].FF/Q REGF\[14\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[7] sky130_fd_sc_hd__ebufn_2
Xfill_7_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[28\].RFW.BIT\[25\].OBUF2 REGF\[28\].RFW.BIT\[25\].FF/Q REGF\[28\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[25] sky130_fd_sc_hd__ebufn_2
XREGF\[20\].RFW.BIT\[27\].OBUF1 REGF\[20\].RFW.BIT\[27\].FF/Q REGF\[20\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[27] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[8\].FF REGF\[27\].RFW.CG\[1\]/GCLK DW[8] VGND VGND VPWR VPWR
+ REGF\[27\].RFW.BIT\[8\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[5\].RFW.BIT\[17\].OBUF1 REGF\[5\].RFW.BIT\[17\].FF/Q REGF\[5\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[17] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.BIT\[6\].OBUF2 REGF\[4\].RFW.BIT\[6\].FF/Q REGF\[4\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[6] sky130_fd_sc_hd__ebufn_2
XREGF\[6\].RFW.BIT\[30\].OBUF1 REGF\[6\].RFW.BIT\[30\].FF/Q REGF\[6\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[30] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.BIT\[23\].OBUF1 REGF\[18\].RFW.BIT\[23\].FF/Q REGF\[18\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[23] sky130_fd_sc_hd__ebufn_2
Xtap_24_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.BIT\[3\].OBUF1 REGF\[18\].RFW.BIT\[3\].FF/Q REGF\[18\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[3] sky130_fd_sc_hd__ebufn_2
Xtap_0_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[23\].RFW.BIT\[12\].OBUF1 REGF\[23\].RFW.BIT\[12\].FF/Q REGF\[23\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[12] sky130_fd_sc_hd__ebufn_2
Xfill_26_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_26_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_26_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[8\].RFW.CG\[1\] CLK REGF\[8\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[8\].RFW.CG\[1\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_42_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_42_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_42_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[8\].RFW.BIT\[2\].OBUF1 REGF\[8\].RFW.BIT\[2\].FF/Q REGF\[8\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[2] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[28\].OBUF2 REGF\[24\].RFW.BIT\[28\].FF/Q REGF\[24\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[28] sky130_fd_sc_hd__ebufn_2
Xtap_50_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_43_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[11\].RFW.BIT\[1\].OBUF1 REGF\[11\].RFW.BIT\[1\].FF/Q REGF\[11\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[1] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[7\].OBUF2 REGF\[16\].RFW.BIT\[7\].FF/Q REGF\[16\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[7] sky130_fd_sc_hd__ebufn_2
XREGF\[30\].RFW.BIT\[30\].OBUF2 REGF\[30\].RFW.BIT\[30\].FF/Q REGF\[30\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[30] sky130_fd_sc_hd__ebufn_2
XREGF\[9\].RFW.BIT\[18\].OBUF2 REGF\[9\].RFW.BIT\[18\].FF/Q REGF\[9\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[18] sky130_fd_sc_hd__ebufn_2
XREGF\[15\].RFW.INV2\[3\] DEC1.D1.AND7/X VGND VGND VPWR VPWR REGF\[15\].RFW.INV2\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[6\].RFW.BIT\[27\].FF REGF\[6\].RFW.CG\[3\]/GCLK DW[27] VGND VGND VPWR VPWR
+ REGF\[6\].RFW.BIT\[27\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[12\].RFW.BIT\[17\].FF REGF\[12\].RFW.CG\[2\]/GCLK DW[17] VGND VGND VPWR VPWR
+ REGF\[12\].RFW.BIT\[17\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[14\].RFW.BIT\[26\].OBUF1 REGF\[14\].RFW.BIT\[26\].FF/Q REGF\[14\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[26] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.BIT\[11\].FF REGF\[18\].RFW.CG\[1\]/GCLK DW[11] VGND VGND VPWR VPWR
+ REGF\[18\].RFW.BIT\[11\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[27\].RFW.BIT\[13\].OBUF2 REGF\[27\].RFW.BIT\[13\].FF/Q REGF\[27\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[13] sky130_fd_sc_hd__ebufn_2
XREGF\[6\].RFW.BIT\[6\].OBUF2 REGF\[6\].RFW.BIT\[6\].FF/Q REGF\[6\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[6] sky130_fd_sc_hd__ebufn_2
XREGF\[1\].RFW.BIT\[0\].OBUF1 REGF\[1\].RFW.BIT\[0\].FF/Q REGF\[1\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[0] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.BIT\[11\].OBUF1 REGF\[17\].RFW.BIT\[11\].FF/Q REGF\[17\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[11] sky130_fd_sc_hd__ebufn_2
XREGF\[8\].RFW.INV1\[0\] DEC0.D1.AND0/Y VGND VGND VPWR VPWR REGF\[8\].RFW.INV1\[0\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_57_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[23\].RFW.BIT\[27\].FF REGF\[23\].RFW.CG\[3\]/GCLK DW[27] VGND VGND VPWR VPWR
+ REGF\[23\].RFW.BIT\[27\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_5_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[29\].RFW.BIT\[21\].FF REGF\[29\].RFW.CG\[2\]/GCLK DW[21] VGND VGND VPWR VPWR
+ REGF\[29\].RFW.BIT\[21\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[18\].RFW.BIT\[27\].OBUF2 REGF\[18\].RFW.BIT\[27\].FF/Q REGF\[18\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[27] sky130_fd_sc_hd__ebufn_2
XREGF\[13\].RFW.BIT\[1\].OBUF1 REGF\[13\].RFW.BIT\[1\].FF/Q REGF\[13\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[1] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.BIT\[7\].OBUF2 REGF\[18\].RFW.BIT\[7\].FF/Q REGF\[18\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[7] sky130_fd_sc_hd__ebufn_2
Xfill_12_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_12_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[10\].RFW.BIT\[29\].OBUF1 REGF\[10\].RFW.BIT\[29\].FF/Q REGF\[10\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[29] sky130_fd_sc_hd__ebufn_2
XREGF\[23\].RFW.BIT\[16\].OBUF2 REGF\[23\].RFW.BIT\[16\].FF/Q REGF\[23\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[16] sky130_fd_sc_hd__ebufn_2
Xtap_22_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[8\].RFW.BIT\[6\].OBUF2 REGF\[8\].RFW.BIT\[6\].FF/Q REGF\[8\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[6] sky130_fd_sc_hd__ebufn_2
XREGF\[1\].RFW.BIT\[21\].OBUF1 REGF\[1\].RFW.BIT\[21\].FF/Q REGF\[1\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[21] sky130_fd_sc_hd__ebufn_2
Xtap_15_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_37_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_37_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XREGF\[3\].RFW.BIT\[0\].OBUF1 REGF\[3\].RFW.BIT\[0\].FF/Q REGF\[3\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[0] sky130_fd_sc_hd__ebufn_2
XREGF\[13\].RFW.BIT\[14\].OBUF1 REGF\[13\].RFW.BIT\[14\].FF/Q REGF\[13\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[14] sky130_fd_sc_hd__ebufn_2
Xtap_8_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_37_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_37_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_37_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[3\].RFW.BIT\[12\].FF REGF\[3\].RFW.CG\[1\]/GCLK DW[12] VGND VGND VPWR VPWR
+ REGF\[3\].RFW.BIT\[12\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_53_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_53_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_53_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_53_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[11\].RFW.BIT\[5\].OBUF2 REGF\[11\].RFW.BIT\[5\].FF/Q REGF\[11\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[5] sky130_fd_sc_hd__ebufn_2
Xfill_53_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC2.D0.AND0 DEC2.D0.AND7/A DEC2.D0.AND7/B DEC2.D0.AND7/C DEC2.D0.AND7/D VGND VGND
+ VPWR VPWR DEC2.D0.AND0/Y sky130_fd_sc_hd__nor4b_2
Xfill_9_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_9_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_9_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[1\].RFW.BIT\[4\].OBUF2 REGF\[1\].RFW.BIT\[4\].FF/Q REGF\[1\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[4] sky130_fd_sc_hd__ebufn_2
Xfill_50_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_43_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_36_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[5\].RFW.BIT\[22\].OBUF2 REGF\[5\].RFW.BIT\[22\].FF/Q REGF\[5\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[22] sky130_fd_sc_hd__ebufn_2
XREGF\[15\].RFW.BIT\[1\].OBUF1 REGF\[15\].RFW.BIT\[1\].FF/Q REGF\[15\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[1] sky130_fd_sc_hd__ebufn_2
Xfill_29_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[17\].RFW.BIT\[15\].OBUF2 REGF\[17\].RFW.BIT\[15\].FF/Q REGF\[17\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[15] sky130_fd_sc_hd__ebufn_2
XREGF\[20\].RFW.BIT\[12\].FF REGF\[20\].RFW.CG\[1\]/GCLK DW[12] VGND VGND VPWR VPWR
+ REGF\[20\].RFW.BIT\[12\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[10\].RFW.BIT\[30\].OBUF1 REGF\[10\].RFW.BIT\[30\].FF/Q REGF\[10\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[30] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[0\].OBUF1 REGF\[5\].RFW.BIT\[0\].FF/Q REGF\[5\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[0] sky130_fd_sc_hd__ebufn_2
Xfill_62_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[13\].RFW.BIT\[5\].OBUF2 REGF\[13\].RFW.BIT\[5\].FF/Q REGF\[13\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[5] sky130_fd_sc_hd__ebufn_2
XREGF\[2\].RFW.INV2\[1\] DEC1.D0.AND2/X VGND VGND VPWR VPWR REGF\[2\].RFW.INV2\[1\]/Y
+ sky130_fd_sc_hd__inv_4
XDEC1.D1.AND2 DEC1.D1.AND7/C DEC1.D1.AND7/A DEC1.D1.AND7/B DEC1.D1.AND7/D VGND VGND
+ VPWR VPWR DEC1.D1.AND2/X sky130_fd_sc_hd__and4bb_2
XREGF\[19\].RFW.BIT\[17\].FF REGF\[19\].RFW.CG\[2\]/GCLK DW[17] VGND VGND VPWR VPWR
+ REGF\[19\].RFW.BIT\[17\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[31\].RFW.BIT\[22\].FF REGF\[31\].RFW.CG\[2\]/GCLK DW[22] VGND VGND VPWR VPWR
+ REGF\[31\].RFW.BIT\[22\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_23_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_23_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_23_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xtap_6_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[1\].RFW.BIT\[25\].OBUF2 REGF\[1\].RFW.BIT\[25\].FF/Q REGF\[1\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[25] sky130_fd_sc_hd__ebufn_2
Xfill_23_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.BIT\[4\].OBUF2 REGF\[3\].RFW.BIT\[4\].FF/Q REGF\[3\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[4] sky130_fd_sc_hd__ebufn_2
XREGF\[14\].RFW.BIT\[31\].OBUF2 REGF\[14\].RFW.BIT\[31\].FF/Q REGF\[14\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[31] sky130_fd_sc_hd__ebufn_2
XREGF\[13\].RFW.BIT\[18\].OBUF2 REGF\[13\].RFW.BIT\[18\].FF/Q REGF\[13\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[18] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.BIT\[1\].OBUF1 REGF\[17\].RFW.BIT\[1\].FF/Q REGF\[17\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[1] sky130_fd_sc_hd__ebufn_2
Xtap_20_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_48_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_48_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_48_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgenblk1.RFW0.BIT\[5\].OBUF1 genblk1.RFW0.TIE\[0\]/LO genblk1.RFW0.INV1\[0\]/Y VGND
+ VGND VPWR VPWR DA[5] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.BIT\[10\].OBUF2 REGF\[4\].RFW.BIT\[10\].FF/Q REGF\[4\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[10] sky130_fd_sc_hd__ebufn_2
XREGF\[11\].RFW.BIT\[1\].FF REGF\[11\].RFW.CG\[0\]/GCLK DW[1] VGND VGND VPWR VPWR
+ REGF\[11\].RFW.BIT\[1\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_6_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[29\].RFW.BIT\[28\].OBUF1 REGF\[29\].RFW.BIT\[28\].FF/Q REGF\[29\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[28] sky130_fd_sc_hd__ebufn_2
XREGF\[7\].RFW.BIT\[0\].OBUF1 REGF\[7\].RFW.BIT\[0\].FF/Q REGF\[7\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[0] sky130_fd_sc_hd__ebufn_2
Xfill_13_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC0.D2.AND4 DEC0.D2.AND7/A DEC0.D2.AND7/B DEC0.D2.AND7/C DEC0.D2.AND7/D VGND VGND
+ VPWR VPWR DEC0.D2.AND4/X sky130_fd_sc_hd__and4bb_2
XREGF\[10\].RFW.BIT\[3\].FF REGF\[10\].RFW.CG\[0\]/GCLK DW[3] VGND VGND VPWR VPWR
+ REGF\[10\].RFW.BIT\[3\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[15\].RFW.BIT\[5\].OBUF2 REGF\[15\].RFW.BIT\[5\].FF/Q REGF\[15\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[5] sky130_fd_sc_hd__ebufn_2
Xfill_41_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_34_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[5\].RFW.BIT\[4\].OBUF2 REGF\[5\].RFW.BIT\[4\].FF/Q REGF\[5\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[4] sky130_fd_sc_hd__ebufn_2
Xfill_27_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[4\].RFW.BIT\[18\].FF REGF\[4\].RFW.CG\[2\]/GCLK DW[18] VGND VGND VPWR VPWR
+ REGF\[4\].RFW.BIT\[18\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_1_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XREGF\[19\].RFW.BIT\[1\].OBUF1 REGF\[19\].RFW.BIT\[1\].FF/Q REGF\[19\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[1] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[1\].FF REGF\[24\].RFW.CG\[0\]/GCLK DW[1] VGND VGND VPWR VPWR
+ REGF\[24\].RFW.BIT\[1\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_18_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_18_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[9\].RFW.BIT\[0\].OBUF1 REGF\[9\].RFW.BIT\[0\].FF/Q REGF\[9\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[0] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.BIT\[18\].FF REGF\[21\].RFW.CG\[2\]/GCLK DW[18] VGND VGND VPWR VPWR
+ REGF\[21\].RFW.BIT\[18\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[28\].RFW.BIT\[16\].OBUF1 REGF\[28\].RFW.BIT\[16\].FF/Q REGF\[28\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[16] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.BIT\[5\].OBUF2 REGF\[17\].RFW.BIT\[5\].FF/Q REGF\[17\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[5] sky130_fd_sc_hd__ebufn_2
Xfill_34_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_34_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xgenblk1.RFW0.BIT\[9\].OBUF2 genblk1.RFW0.TIE\[5\]/LO genblk1.RFW0.INV2\[1\]/Y VGND
+ VGND VPWR VPWR DB[9] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.INV2\[0\] DEC1.D2.AND1/X VGND VGND VPWR VPWR REGF\[17\].RFW.INV2\[0\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[27\].RFW.BIT\[12\].FF REGF\[27\].RFW.CG\[1\]/GCLK DW[12] VGND VGND VPWR VPWR
+ REGF\[27\].RFW.BIT\[12\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_50_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_50_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[23\].RFW.BIT\[3\].FF REGF\[23\].RFW.CG\[0\]/GCLK DW[3] VGND VGND VPWR VPWR
+ REGF\[23\].RFW.BIT\[3\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_50_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_59_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_59_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_59_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_59_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_6_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_59_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[7\].RFW.BIT\[4\].OBUF2 REGF\[7\].RFW.BIT\[4\].FF/Q REGF\[7\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[4] sky130_fd_sc_hd__ebufn_2
XREGF\[10\].RFW.BIT\[3\].OBUF2 REGF\[10\].RFW.BIT\[3\].FF/Q REGF\[10\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[3] sky130_fd_sc_hd__ebufn_2
Xfill_13_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[16\].RFW.BIT\[25\].FF REGF\[16\].RFW.CG\[3\]/GCLK DW[25] VGND VGND VPWR VPWR
+ REGF\[16\].RFW.BIT\[25\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[22\].RFW.BIT\[5\].FF REGF\[22\].RFW.CG\[0\]/GCLK DW[5] VGND VGND VPWR VPWR
+ REGF\[22\].RFW.BIT\[5\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[24\].RFW.BIT\[19\].OBUF1 REGF\[24\].RFW.BIT\[19\].FF/Q REGF\[24\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[19] sky130_fd_sc_hd__ebufn_2
XREGF\[8\].RFW.BIT\[0\].FF REGF\[8\].RFW.CG\[0\]/GCLK DW[0] VGND VGND VPWR VPWR REGF\[8\].RFW.BIT\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[30\].RFW.BIT\[21\].OBUF1 REGF\[30\].RFW.BIT\[21\].FF/Q REGF\[30\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[21] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.BIT\[7\].FF REGF\[21\].RFW.CG\[0\]/GCLK DW[7] VGND VGND VPWR VPWR
+ REGF\[21\].RFW.BIT\[7\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[19\].RFW.BIT\[5\].OBUF2 REGF\[19\].RFW.BIT\[5\].FF/Q REGF\[19\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[5] sky130_fd_sc_hd__ebufn_2
Xfill_32_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[13\].RFW.INV1\[1\] DEC0.D1.AND5/X VGND VGND VPWR VPWR REGF\[13\].RFW.INV1\[1\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_25_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[21\].RFW.BIT\[8\].OBUF1 REGF\[21\].RFW.BIT\[8\].FF/Q REGF\[21\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[8] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.INV1\[2\] DEC0.D3.AND5/X VGND VGND VPWR VPWR REGF\[29\].RFW.INV1\[2\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[7\].RFW.BIT\[2\].FF REGF\[7\].RFW.CG\[0\]/GCLK DW[2] VGND VGND VPWR VPWR REGF\[7\].RFW.BIT\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[9\].RFW.BIT\[4\].OBUF2 REGF\[9\].RFW.BIT\[4\].FF/Q REGF\[9\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[4] sky130_fd_sc_hd__ebufn_2
Xtap_54_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_20_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[9\].FF REGF\[20\].RFW.CG\[1\]/GCLK DW[9] VGND VGND VPWR VPWR
+ REGF\[20\].RFW.BIT\[9\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_20_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.BIT\[3\].OBUF2 REGF\[12\].RFW.BIT\[3\].FF/Q REGF\[12\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[3] sky130_fd_sc_hd__ebufn_2
Xfill_29_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_29_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_29_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_29_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_29_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_45_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.BIT\[25\].OBUF1 REGF\[6\].RFW.BIT\[25\].FF/Q REGF\[6\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[25] sky130_fd_sc_hd__ebufn_2
XREGF\[6\].RFW.BIT\[4\].FF REGF\[6\].RFW.CG\[0\]/GCLK DW[4] VGND VGND VPWR VPWR REGF\[6\].RFW.BIT\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[1\].RFW.BIT\[26\].FF REGF\[1\].RFW.CG\[3\]/GCLK DW[26] VGND VGND VPWR VPWR
+ REGF\[1\].RFW.BIT\[26\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_45_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_45_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_45_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_45_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[18\].RFW.BIT\[18\].OBUF1 REGF\[18\].RFW.BIT\[18\].FF/Q REGF\[18\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[18] sky130_fd_sc_hd__ebufn_2
Xfill_61_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_61_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_61_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[7\].RFW.BIT\[20\].FF REGF\[7\].RFW.CG\[2\]/GCLK DW[20] VGND VGND VPWR VPWR
+ REGF\[7\].RFW.BIT\[20\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[13\].RFW.BIT\[10\].FF REGF\[13\].RFW.CG\[1\]/GCLK DW[10] VGND VGND VPWR VPWR
+ REGF\[13\].RFW.BIT\[10\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[19\].RFW.BIT\[31\].OBUF1 REGF\[19\].RFW.BIT\[31\].FF/Q REGF\[19\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[31] sky130_fd_sc_hd__ebufn_2
Xfill_61_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_61_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[2\].RFW.BIT\[2\].OBUF2 REGF\[2\].RFW.BIT\[2\].FF/Q REGF\[2\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[2] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[20\].OBUF1 REGF\[24\].RFW.BIT\[20\].FF/Q REGF\[24\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[20] sky130_fd_sc_hd__ebufn_2
XREGF\[9\].RFW.BIT\[10\].OBUF1 REGF\[9\].RFW.BIT\[10\].FF/Q REGF\[9\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[10] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[6\].FF REGF\[5\].RFW.CG\[0\]/GCLK DW[6] VGND VGND VPWR VPWR REGF\[5\].RFW.BIT\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[5\].RFW.CG\[3\] CLK REGF\[5\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[5\].RFW.CG\[3\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[23\].RFW.BIT\[8\].OBUF1 REGF\[23\].RFW.BIT\[8\].FF/Q REGF\[23\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[8] sky130_fd_sc_hd__ebufn_2
Xfill_11_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_9_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[30\].RFW.BIT\[25\].OBUF2 REGF\[30\].RFW.BIT\[25\].FF/Q REGF\[30\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[25] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.BIT\[18\].FF REGF\[28\].RFW.CG\[2\]/GCLK DW[18] VGND VGND VPWR VPWR
+ REGF\[28\].RFW.BIT\[18\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[24\].RFW.BIT\[20\].FF REGF\[24\].RFW.CG\[2\]/GCLK DW[20] VGND VGND VPWR VPWR
+ REGF\[24\].RFW.BIT\[20\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[4\].RFW.BIT\[8\].FF REGF\[4\].RFW.CG\[1\]/GCLK DW[8] VGND VGND VPWR VPWR REGF\[4\].RFW.BIT\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[2\].RFW.BIT\[28\].OBUF1 REGF\[2\].RFW.BIT\[28\].FF/Q REGF\[2\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[28] sky130_fd_sc_hd__ebufn_2
XREGF\[14\].RFW.BIT\[3\].OBUF2 REGF\[14\].RFW.BIT\[3\].FF/Q REGF\[14\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[3] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.BIT\[21\].OBUF2 REGF\[28\].RFW.BIT\[21\].FF/Q REGF\[28\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[21] sky130_fd_sc_hd__ebufn_2
Xfill_7_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_7_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[23\].OBUF1 REGF\[20\].RFW.BIT\[23\].FF/Q REGF\[20\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[23] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.BIT\[2\].OBUF2 REGF\[4\].RFW.BIT\[2\].FF/Q REGF\[4\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[2] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[13\].OBUF1 REGF\[5\].RFW.BIT\[13\].FF/Q REGF\[5\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[13] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.CG\[0\] CLK REGF\[4\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[4\].RFW.CG\[0\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_15_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_15_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_15_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_31_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_31_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[23\].RFW.INV2\[3\] DEC1.D2.AND7/X VGND VGND VPWR VPWR REGF\[23\].RFW.INV2\[3\]/Y
+ sky130_fd_sc_hd__inv_4
Xtap_52_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_31_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_31_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.BIT\[29\].OBUF2 REGF\[6\].RFW.BIT\[29\].FF/Q REGF\[6\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[29] sky130_fd_sc_hd__ebufn_2
XREGF\[25\].RFW.BIT\[8\].OBUF1 REGF\[25\].RFW.BIT\[8\].FF/Q REGF\[25\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[8] sky130_fd_sc_hd__ebufn_2
Xtap_38_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_56_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_56_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_56_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[24\].RFW.BIT\[24\].OBUF2 REGF\[24\].RFW.BIT\[24\].FF/Q REGF\[24\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[24] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[3\].OBUF2 REGF\[16\].RFW.BIT\[3\].FF/Q REGF\[16\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[3] sky130_fd_sc_hd__ebufn_2
XREGF\[9\].RFW.BIT\[14\].OBUF2 REGF\[9\].RFW.BIT\[14\].FF/Q REGF\[9\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[14] sky130_fd_sc_hd__ebufn_2
XREGF\[1\].RFW.BIT\[16\].OBUF1 REGF\[1\].RFW.BIT\[16\].FF/Q REGF\[1\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[16] sky130_fd_sc_hd__ebufn_2
XREGF\[14\].RFW.BIT\[22\].OBUF1 REGF\[14\].RFW.BIT\[22\].FF/Q REGF\[14\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[22] sky130_fd_sc_hd__ebufn_2
Xfill_21_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.BIT\[2\].OBUF2 REGF\[6\].RFW.BIT\[2\].FF/Q REGF\[6\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[2] sky130_fd_sc_hd__ebufn_2
Xfill_59_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_7_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[8\].RFW.BIT\[26\].FF REGF\[8\].RFW.CG\[3\]/GCLK DW[26] VGND VGND VPWR VPWR
+ REGF\[8\].RFW.BIT\[26\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[14\].RFW.BIT\[16\].FF REGF\[14\].RFW.CG\[2\]/GCLK DW[16] VGND VGND VPWR VPWR
+ REGF\[14\].RFW.BIT\[16\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[19\].RFW.CG\[2\] CLK REGF\[19\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[19\].RFW.CG\[2\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[20\].RFW.BIT\[27\].OBUF2 REGF\[20\].RFW.BIT\[27\].FF/Q REGF\[20\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[27] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[8\].OBUF1 REGF\[27\].RFW.BIT\[8\].FF/Q REGF\[27\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[8] sky130_fd_sc_hd__ebufn_2
XREGF\[30\].RFW.BIT\[19\].FF REGF\[30\].RFW.CG\[2\]/GCLK DW[19] VGND VGND VPWR VPWR
+ REGF\[30\].RFW.BIT\[19\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[6\].RFW.BIT\[30\].OBUF2 REGF\[6\].RFW.BIT\[30\].FF/Q REGF\[6\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[30] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[17\].OBUF2 REGF\[5\].RFW.BIT\[17\].FF/Q REGF\[5\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[17] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.BIT\[23\].OBUF2 REGF\[18\].RFW.BIT\[23\].FF/Q REGF\[18\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[23] sky130_fd_sc_hd__ebufn_2
Xtap_24_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.BIT\[3\].OBUF2 REGF\[18\].RFW.BIT\[3\].FF/Q REGF\[18\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[3] sky130_fd_sc_hd__ebufn_2
XREGF\[10\].RFW.BIT\[25\].OBUF1 REGF\[10\].RFW.BIT\[25\].FF/Q REGF\[10\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[25] sky130_fd_sc_hd__ebufn_2
Xtap_0_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[23\].RFW.BIT\[12\].OBUF2 REGF\[23\].RFW.BIT\[12\].FF/Q REGF\[23\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[12] sky130_fd_sc_hd__ebufn_2
Xfill_26_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_26_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[6\].OBUF1 REGF\[20\].RFW.BIT\[6\].FF/Q REGF\[20\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[6] sky130_fd_sc_hd__ebufn_2
XREGF\[25\].RFW.BIT\[26\].FF REGF\[25\].RFW.CG\[3\]/GCLK DW[26] VGND VGND VPWR VPWR
+ REGF\[25\].RFW.BIT\[26\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_42_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_42_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[8\].RFW.BIT\[2\].OBUF2 REGF\[8\].RFW.BIT\[2\].FF/Q REGF\[8\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[2] sky130_fd_sc_hd__ebufn_2
Xfill_42_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[13\].RFW.BIT\[10\].OBUF1 REGF\[13\].RFW.BIT\[10\].FF/Q REGF\[13\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[10] sky130_fd_sc_hd__ebufn_2
Xtap_50_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_43_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_36_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[11\].RFW.BIT\[1\].OBUF2 REGF\[11\].RFW.BIT\[1\].FF/Q REGF\[11\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[1] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.BIT\[8\].OBUF1 REGF\[29\].RFW.BIT\[8\].FF/Q REGF\[29\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[8] sky130_fd_sc_hd__ebufn_2
XREGF\[14\].RFW.BIT\[26\].OBUF2 REGF\[14\].RFW.BIT\[26\].FF/Q REGF\[14\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[26] sky130_fd_sc_hd__ebufn_2
XREGF\[1\].RFW.BIT\[0\].OBUF2 REGF\[1\].RFW.BIT\[0\].FF/Q REGF\[1\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[0] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[11\].FF REGF\[5\].RFW.CG\[1\]/GCLK DW[11] VGND VGND VPWR VPWR
+ REGF\[5\].RFW.BIT\[11\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[17\].RFW.BIT\[11\].OBUF2 REGF\[17\].RFW.BIT\[11\].FF/Q REGF\[17\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[11] sky130_fd_sc_hd__ebufn_2
Xfill_57_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[22\].RFW.BIT\[6\].OBUF1 REGF\[22\].RFW.BIT\[6\].FF/Q REGF\[22\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[6] sky130_fd_sc_hd__ebufn_2
Xfill_5_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XREGF\[13\].RFW.BIT\[1\].OBUF2 REGF\[13\].RFW.BIT\[1\].FF/Q REGF\[13\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[1] sky130_fd_sc_hd__ebufn_2
Xfill_12_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[10\].RFW.BIT\[29\].OBUF2 REGF\[10\].RFW.BIT\[29\].FF/Q REGF\[10\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[29] sky130_fd_sc_hd__ebufn_2
Xfill_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[22\].RFW.BIT\[11\].FF REGF\[22\].RFW.CG\[1\]/GCLK DW[11] VGND VGND VPWR VPWR
+ REGF\[22\].RFW.BIT\[11\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_22_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[1\].RFW.BIT\[21\].OBUF2 REGF\[1\].RFW.BIT\[21\].FF/Q REGF\[1\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[21] sky130_fd_sc_hd__ebufn_2
Xfill_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[3\].RFW.BIT\[0\].OBUF2 REGF\[3\].RFW.BIT\[0\].FF/Q REGF\[3\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[0] sky130_fd_sc_hd__ebufn_2
XREGF\[13\].RFW.BIT\[14\].OBUF2 REGF\[13\].RFW.BIT\[14\].FF/Q REGF\[13\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[14] sky130_fd_sc_hd__ebufn_2
Xtap_8_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_37_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_37_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_37_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_37_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_53_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_53_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_53_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_53_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_53_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.BIT\[28\].OBUF1 REGF\[31\].RFW.BIT\[28\].FF/Q REGF\[31\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[28] sky130_fd_sc_hd__ebufn_2
XREGF\[11\].RFW.BIT\[24\].FF REGF\[11\].RFW.CG\[3\]/GCLK DW[24] VGND VGND VPWR VPWR
+ REGF\[11\].RFW.BIT\[24\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xgenblk1.RFW0.BIT\[1\].OBUF1 genblk1.RFW0.TIE\[0\]/LO genblk1.RFW0.INV1\[0\]/Y VGND
+ VGND VPWR VPWR DA[1] sky130_fd_sc_hd__ebufn_2
XDEC2.D0.AND1 DEC2.D0.AND7/C DEC2.D0.AND7/B DEC2.D0.AND7/A DEC2.D0.AND7/D VGND VGND
+ VPWR VPWR DEC2.D0.AND1/X sky130_fd_sc_hd__and4bb_2
XDEC2.D1.ABUF\[2\] RW[2] VGND VGND VPWR VPWR DEC2.D1.AND7/C sky130_fd_sc_hd__clkbuf_2
Xfill_9_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_9_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[24\].RFW.BIT\[6\].OBUF1 REGF\[24\].RFW.BIT\[6\].FF/Q REGF\[24\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[6] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.BIT\[24\].OBUF1 REGF\[29\].RFW.BIT\[24\].FF/Q REGF\[29\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[24] sky130_fd_sc_hd__ebufn_2
Xfill_43_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_36_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[15\].RFW.BIT\[1\].OBUF2 REGF\[15\].RFW.BIT\[1\].FF/Q REGF\[15\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[1] sky130_fd_sc_hd__ebufn_2
Xfill_29_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[5\].RFW.INV2\[2\] DEC1.D0.AND5/X VGND VGND VPWR VPWR REGF\[5\].RFW.INV2\[2\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[31\].RFW.BIT\[0\].FF REGF\[31\].RFW.CG\[0\]/GCLK DW[0] VGND VGND VPWR VPWR
+ REGF\[31\].RFW.BIT\[0\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[10\].RFW.BIT\[30\].OBUF2 REGF\[10\].RFW.BIT\[30\].FF/Q REGF\[10\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[30] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[0\].OBUF2 REGF\[5\].RFW.BIT\[0\].FF/Q REGF\[5\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[0] sky130_fd_sc_hd__ebufn_2
Xfill_62_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_55_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC1.D1.AND3 DEC1.D1.AND7/C DEC1.D1.AND7/B DEC1.D1.AND7/A DEC1.D1.AND7/D VGND VGND
+ VPWR VPWR DEC1.D1.AND3/X sky130_fd_sc_hd__and4b_2
XREGF\[30\].RFW.BIT\[2\].FF REGF\[30\].RFW.CG\[0\]/GCLK DW[2] VGND VGND VPWR VPWR
+ REGF\[30\].RFW.BIT\[2\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[1\].RFW.BIT\[1\].FF REGF\[1\].RFW.CG\[0\]/GCLK DW[1] VGND VGND VPWR VPWR REGF\[1\].RFW.BIT\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[25\].RFW.BIT\[27\].OBUF1 REGF\[25\].RFW.BIT\[27\].FF/Q REGF\[25\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[27] sky130_fd_sc_hd__ebufn_2
XREGF\[25\].RFW.INV2\[0\] DEC1.D3.AND1/X VGND VGND VPWR VPWR REGF\[25\].RFW.INV2\[0\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[30\].RFW.BIT\[16\].OBUF1 REGF\[30\].RFW.BIT\[16\].FF/Q REGF\[30\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[16] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[6\].OBUF1 REGF\[26\].RFW.BIT\[6\].FF/Q REGF\[26\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[6] sky130_fd_sc_hd__ebufn_2
Xfill_23_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_23_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xtap_6_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_23_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.BIT\[17\].FF REGF\[6\].RFW.CG\[2\]/GCLK DW[17] VGND VGND VPWR VPWR
+ REGF\[6\].RFW.BIT\[17\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[28\].RFW.BIT\[12\].OBUF1 REGF\[28\].RFW.BIT\[12\].FF/Q REGF\[28\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[12] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.BIT\[1\].OBUF2 REGF\[17\].RFW.BIT\[1\].FF/Q REGF\[17\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[1] sky130_fd_sc_hd__ebufn_2
Xtap_20_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_48_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_48_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgenblk1.RFW0.BIT\[5\].OBUF2 genblk1.RFW0.TIE\[4\]/LO genblk1.RFW0.INV2\[0\]/Y VGND
+ VGND VPWR VPWR DB[5] sky130_fd_sc_hd__ebufn_2
Xfill_48_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[1\].RFW.INV1\[3\] DEC0.D0.AND1/X VGND VGND VPWR VPWR REGF\[1\].RFW.INV1\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[29\].RFW.BIT\[28\].OBUF2 REGF\[29\].RFW.BIT\[28\].FF/Q REGF\[29\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[28] sky130_fd_sc_hd__ebufn_2
XREGF\[7\].RFW.BIT\[0\].OBUF2 REGF\[7\].RFW.BIT\[0\].FF/Q REGF\[7\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[0] sky130_fd_sc_hd__ebufn_2
Xfill_13_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_13_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDEC0.D2.AND5 DEC0.D2.AND7/B DEC0.D2.AND7/A DEC0.D2.AND7/C DEC0.D2.AND7/D VGND VGND
+ VPWR VPWR DEC0.D2.AND5/X sky130_fd_sc_hd__and4b_2
XREGF\[23\].RFW.BIT\[17\].FF REGF\[23\].RFW.CG\[2\]/GCLK DW[17] VGND VGND VPWR VPWR
+ REGF\[23\].RFW.BIT\[17\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[29\].RFW.BIT\[11\].FF REGF\[29\].RFW.CG\[1\]/GCLK DW[11] VGND VGND VPWR VPWR
+ REGF\[29\].RFW.BIT\[11\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[19\].RFW.BIT\[26\].OBUF1 REGF\[19\].RFW.BIT\[26\].FF/Q REGF\[19\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[26] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.INV1\[1\] DEC0.D2.AND5/X VGND VGND VPWR VPWR REGF\[21\].RFW.INV1\[1\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_41_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[28\].RFW.BIT\[6\].OBUF1 REGF\[28\].RFW.BIT\[6\].FF/Q REGF\[28\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[6] sky130_fd_sc_hd__ebufn_2
Xfill_34_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[24\].RFW.BIT\[15\].OBUF1 REGF\[24\].RFW.BIT\[15\].FF/Q REGF\[24\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[15] sky130_fd_sc_hd__ebufn_2
Xfill_27_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[19\].RFW.BIT\[1\].OBUF2 REGF\[19\].RFW.BIT\[1\].FF/Q REGF\[19\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[1] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.BIT\[24\].FF REGF\[18\].RFW.CG\[3\]/GCLK DW[24] VGND VGND VPWR VPWR
+ REGF\[18\].RFW.BIT\[24\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[21\].RFW.BIT\[4\].OBUF1 REGF\[21\].RFW.BIT\[4\].FF/Q REGF\[21\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[4] sky130_fd_sc_hd__ebufn_2
Xfill_18_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[9\].RFW.BIT\[0\].OBUF2 REGF\[9\].RFW.BIT\[0\].FF/Q REGF\[9\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[0] sky130_fd_sc_hd__ebufn_2
Xfill_18_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[15\].RFW.BIT\[29\].OBUF1 REGF\[15\].RFW.BIT\[29\].FF/Q REGF\[15\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[29] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.BIT\[16\].OBUF2 REGF\[28\].RFW.BIT\[16\].FF/Q REGF\[28\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[16] sky130_fd_sc_hd__ebufn_2
Xfill_34_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[20\].RFW.BIT\[18\].OBUF1 REGF\[20\].RFW.BIT\[18\].FF/Q REGF\[20\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[18] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.BIT\[31\].OBUF1 REGF\[21\].RFW.BIT\[31\].FF/Q REGF\[21\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[31] sky130_fd_sc_hd__ebufn_2
Xfill_50_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_50_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_50_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[6\].RFW.BIT\[21\].OBUF1 REGF\[6\].RFW.BIT\[21\].FF/Q REGF\[6\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[21] sky130_fd_sc_hd__ebufn_2
Xfill_59_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_59_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_59_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_6_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_59_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_59_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[1\].RFW.CG\[2\] CLK REGF\[1\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[1\].RFW.CG\[2\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[18\].RFW.BIT\[14\].OBUF1 REGF\[18\].RFW.BIT\[14\].FF/Q REGF\[18\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[14] sky130_fd_sc_hd__ebufn_2
XREGF\[23\].RFW.BIT\[4\].OBUF1 REGF\[23\].RFW.BIT\[4\].FF/Q REGF\[23\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[4] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[19\].OBUF2 REGF\[24\].RFW.BIT\[19\].FF/Q REGF\[24\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[19] sky130_fd_sc_hd__ebufn_2
XREGF\[3\].RFW.BIT\[25\].FF REGF\[3\].RFW.CG\[3\]/GCLK DW[25] VGND VGND VPWR VPWR
+ REGF\[3\].RFW.BIT\[25\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[27\].RFW.CG\[1\] CLK REGF\[27\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[27\].RFW.CG\[1\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[16\].RFW.INV1\[2\] DEC0.D2.AND0/Y VGND VGND VPWR VPWR REGF\[16\].RFW.INV1\[2\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[30\].RFW.BIT\[21\].OBUF2 REGF\[30\].RFW.BIT\[21\].FF/Q REGF\[30\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[21] sky130_fd_sc_hd__ebufn_2
XREGF\[31\].RFW.BIT\[12\].FF REGF\[31\].RFW.CG\[1\]/GCLK DW[12] VGND VGND VPWR VPWR
+ REGF\[31\].RFW.BIT\[12\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[2\].RFW.BIT\[24\].OBUF1 REGF\[2\].RFW.BIT\[24\].FF/Q REGF\[2\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[24] sky130_fd_sc_hd__ebufn_2
Xfill_32_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[14\].RFW.BIT\[17\].OBUF1 REGF\[14\].RFW.BIT\[17\].FF/Q REGF\[14\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[17] sky130_fd_sc_hd__ebufn_2
XREGF\[15\].RFW.BIT\[30\].OBUF1 REGF\[15\].RFW.BIT\[30\].FF/Q REGF\[15\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[30] sky130_fd_sc_hd__ebufn_2
Xfill_25_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_18_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.INV2\[3\] DEC1.D3.AND7/X VGND VGND VPWR VPWR REGF\[31\].RFW.INV2\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[21\].RFW.BIT\[8\].OBUF2 REGF\[21\].RFW.BIT\[8\].FF/Q REGF\[21\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[8] sky130_fd_sc_hd__ebufn_2
Xtap_54_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[25\].FF REGF\[20\].RFW.CG\[3\]/GCLK DW[25] VGND VGND VPWR VPWR
+ REGF\[20\].RFW.BIT\[25\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_20_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_29_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_29_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_29_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_29_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_45_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_45_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_45_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[6\].RFW.BIT\[25\].OBUF2 REGF\[6\].RFW.BIT\[25\].FF/Q REGF\[6\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[25] sky130_fd_sc_hd__ebufn_2
XREGF\[25\].RFW.BIT\[4\].OBUF1 REGF\[25\].RFW.BIT\[4\].FF/Q REGF\[25\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[4] sky130_fd_sc_hd__ebufn_2
Xfill_45_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.BIT\[18\].OBUF2 REGF\[18\].RFW.BIT\[18\].FF/Q REGF\[18\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[18] sky130_fd_sc_hd__ebufn_2
Xfill_61_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_61_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[19\].RFW.BIT\[31\].OBUF2 REGF\[19\].RFW.BIT\[31\].FF/Q REGF\[19\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[31] sky130_fd_sc_hd__ebufn_2
Xfill_61_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_61_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_61_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[24\].RFW.BIT\[20\].OBUF2 REGF\[24\].RFW.BIT\[20\].FF/Q REGF\[24\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[20] sky130_fd_sc_hd__ebufn_2
XREGF\[9\].RFW.BIT\[10\].OBUF2 REGF\[9\].RFW.BIT\[10\].FF/Q REGF\[9\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[10] sky130_fd_sc_hd__ebufn_2
XREGF\[1\].RFW.BIT\[12\].OBUF1 REGF\[1\].RFW.BIT\[12\].FF/Q REGF\[1\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[12] sky130_fd_sc_hd__ebufn_2
XREGF\[23\].RFW.BIT\[8\].OBUF2 REGF\[23\].RFW.BIT\[8\].FF/Q REGF\[23\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[8] sky130_fd_sc_hd__ebufn_2
Xfill_19_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_11_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_9_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[15\].RFW.CG\[1\] CLK REGF\[15\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[15\].RFW.CG\[1\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[2\].RFW.BIT\[28\].OBUF2 REGF\[2\].RFW.BIT\[28\].FF/Q REGF\[2\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[28] sky130_fd_sc_hd__ebufn_2
Xfill_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_7_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[10\].RFW.INV2\[3\] DEC1.D1.AND2/X VGND VGND VPWR VPWR REGF\[10\].RFW.INV2\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[20\].RFW.BIT\[23\].OBUF2 REGF\[20\].RFW.BIT\[23\].FF/Q REGF\[20\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[23] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[4\].OBUF1 REGF\[27\].RFW.BIT\[4\].FF/Q REGF\[27\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[4] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[13\].OBUF2 REGF\[5\].RFW.BIT\[13\].FF/Q REGF\[5\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[13] sky130_fd_sc_hd__ebufn_2
Xfill_15_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_15_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[10\].RFW.BIT\[21\].OBUF1 REGF\[10\].RFW.BIT\[21\].FF/Q REGF\[10\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[21] sky130_fd_sc_hd__ebufn_2
Xfill_31_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_52_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_31_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_31_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[16\].RFW.BIT\[15\].FF REGF\[16\].RFW.CG\[1\]/GCLK DW[15] VGND VGND VPWR VPWR
+ REGF\[16\].RFW.BIT\[15\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[25\].RFW.BIT\[8\].OBUF2 REGF\[25\].RFW.BIT\[8\].FF/Q REGF\[25\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[8] sky130_fd_sc_hd__ebufn_2
Xtap_38_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[2\].OBUF1 REGF\[20\].RFW.BIT\[2\].FF/Q REGF\[20\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[2] sky130_fd_sc_hd__ebufn_2
XREGF\[3\].RFW.INV1\[0\] DEC0.D0.AND3/X VGND VGND VPWR VPWR REGF\[3\].RFW.INV1\[0\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_56_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_56_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_56_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[1\].RFW.BIT\[16\].OBUF2 REGF\[1\].RFW.BIT\[16\].FF/Q REGF\[1\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[16] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.BIT\[4\].OBUF1 REGF\[29\].RFW.BIT\[4\].FF/Q REGF\[29\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[4] sky130_fd_sc_hd__ebufn_2
XREGF\[14\].RFW.BIT\[22\].OBUF2 REGF\[14\].RFW.BIT\[22\].FF/Q REGF\[14\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[22] sky130_fd_sc_hd__ebufn_2
Xfill_21_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[27\].RFW.BIT\[25\].FF REGF\[27\].RFW.CG\[3\]/GCLK DW[25] VGND VGND VPWR VPWR
+ REGF\[27\].RFW.BIT\[25\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_59_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgenblk1.RFW0.INV1\[3\] DEC0.D0.AND0/Y VGND VGND VPWR VPWR genblk1.RFW0.INV1\[3\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_7_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[29\].RFW.BIT\[19\].OBUF1 REGF\[29\].RFW.BIT\[19\].FF/Q REGF\[29\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[19] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[8\].OBUF2 REGF\[27\].RFW.BIT\[8\].FF/Q REGF\[27\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[8] sky130_fd_sc_hd__ebufn_2
XREGF\[22\].RFW.BIT\[2\].OBUF1 REGF\[22\].RFW.BIT\[2\].FF/Q REGF\[22\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[2] sky130_fd_sc_hd__ebufn_2
XREGF\[1\].RFW.BIT\[16\].FF REGF\[1\].RFW.CG\[2\]/GCLK DW[16] VGND VGND VPWR VPWR
+ REGF\[1\].RFW.BIT\[16\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[7\].RFW.BIT\[10\].FF REGF\[7\].RFW.CG\[1\]/GCLK DW[10] VGND VGND VPWR VPWR
+ REGF\[7\].RFW.BIT\[10\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[10\].RFW.BIT\[25\].OBUF2 REGF\[10\].RFW.BIT\[25\].FF/Q REGF\[10\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[25] sky130_fd_sc_hd__ebufn_2
Xtap_0_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_26_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_26_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[20\].RFW.BIT\[6\].OBUF2 REGF\[20\].RFW.BIT\[6\].FF/Q REGF\[20\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[6] sky130_fd_sc_hd__ebufn_2
Xfill_42_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_42_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_42_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[13\].RFW.BIT\[10\].OBUF2 REGF\[13\].RFW.BIT\[10\].FF/Q REGF\[13\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[10] sky130_fd_sc_hd__ebufn_2
Xtap_50_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_43_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_36_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.BIT\[24\].OBUF1 REGF\[31\].RFW.BIT\[24\].FF/Q REGF\[31\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[24] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[10\].FF REGF\[24\].RFW.CG\[1\]/GCLK DW[10] VGND VGND VPWR VPWR
+ REGF\[24\].RFW.BIT\[10\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[29\].RFW.BIT\[8\].OBUF2 REGF\[29\].RFW.BIT\[8\].FF/Q REGF\[29\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[8] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[2\].OBUF1 REGF\[24\].RFW.BIT\[2\].FF/Q REGF\[24\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[2] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.BIT\[20\].OBUF1 REGF\[29\].RFW.BIT\[20\].FF/Q REGF\[29\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[20] sky130_fd_sc_hd__ebufn_2
XREGF\[13\].RFW.BIT\[23\].FF REGF\[13\].RFW.CG\[2\]/GCLK DW[23] VGND VGND VPWR VPWR
+ REGF\[13\].RFW.BIT\[23\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xgenblk1.RFW0.TIE\[0\] VGND VGND VPWR VPWR genblk1.RFW0.TIE\[0\]/HI genblk1.RFW0.TIE\[0\]/LO
+ sky130_fd_sc_hd__conb_1
Xfill_57_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[22\].RFW.BIT\[6\].OBUF2 REGF\[22\].RFW.BIT\[6\].FF/Q REGF\[22\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[6] sky130_fd_sc_hd__ebufn_2
Xfill_4_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_5_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[7\].RFW.BIT\[28\].OBUF1 REGF\[7\].RFW.BIT\[28\].FF/Q REGF\[7\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[28] sky130_fd_sc_hd__ebufn_2
Xfill_12_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[25\].RFW.BIT\[23\].OBUF1 REGF\[25\].RFW.BIT\[23\].FF/Q REGF\[25\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[23] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[2\].OBUF1 REGF\[26\].RFW.BIT\[2\].FF/Q REGF\[26\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[2] sky130_fd_sc_hd__ebufn_2
XREGF\[30\].RFW.BIT\[12\].OBUF1 REGF\[30\].RFW.BIT\[12\].FF/Q REGF\[30\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[12] sky130_fd_sc_hd__ebufn_2
Xtap_22_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_37_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_37_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_37_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_53_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_53_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_53_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_53_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_53_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[31\].RFW.BIT\[28\].OBUF2 REGF\[31\].RFW.BIT\[28\].FF/Q REGF\[31\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[28] sky130_fd_sc_hd__ebufn_2
XDEC2.D0.AND2 DEC2.D0.AND7/C DEC2.D0.AND7/A DEC2.D0.AND7/B DEC2.D0.AND7/D VGND VGND
+ VPWR VPWR DEC2.D0.AND2/X sky130_fd_sc_hd__and4bb_2
Xgenblk1.RFW0.BIT\[1\].OBUF2 genblk1.RFW0.TIE\[4\]/LO genblk1.RFW0.INV2\[0\]/Y VGND
+ VGND VPWR VPWR DB[1] sky130_fd_sc_hd__ebufn_2
Xfill_9_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[24\].RFW.BIT\[6\].OBUF2 REGF\[24\].RFW.BIT\[6\].FF/Q REGF\[24\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[6] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.BIT\[24\].OBUF2 REGF\[29\].RFW.BIT\[24\].FF/Q REGF\[29\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[24] sky130_fd_sc_hd__ebufn_2
XREGF\[8\].RFW.INV2\[3\] DEC1.D1.AND0/Y VGND VGND VPWR VPWR REGF\[8\].RFW.INV2\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[8\].RFW.BIT\[16\].FF REGF\[8\].RFW.CG\[2\]/GCLK DW[16] VGND VGND VPWR VPWR
+ REGF\[8\].RFW.BIT\[16\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[21\].RFW.BIT\[26\].OBUF1 REGF\[21\].RFW.BIT\[26\].FF/Q REGF\[21\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[26] sky130_fd_sc_hd__ebufn_2
Xfill_36_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_27_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_29_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[6\].RFW.BIT\[16\].OBUF1 REGF\[6\].RFW.BIT\[16\].FF/Q REGF\[6\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[16] sky130_fd_sc_hd__ebufn_2
XREGF\[12\].RFW.INV2\[0\] DEC1.D1.AND4/X VGND VGND VPWR VPWR REGF\[12\].RFW.INV2\[0\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[19\].RFW.BIT\[22\].OBUF1 REGF\[19\].RFW.BIT\[22\].FF/Q REGF\[19\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[22] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.BIT\[2\].OBUF1 REGF\[28\].RFW.BIT\[2\].FF/Q REGF\[28\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[2] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[11\].OBUF1 REGF\[24\].RFW.BIT\[11\].FF/Q REGF\[24\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[11] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.INV2\[1\] DEC1.D3.AND4/X VGND VGND VPWR VPWR REGF\[28\].RFW.INV2\[1\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_62_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_55_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[19\].RFW.BIT\[1\].FF REGF\[19\].RFW.CG\[0\]/GCLK DW[1] VGND VGND VPWR VPWR
+ REGF\[19\].RFW.BIT\[1\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[25\].RFW.BIT\[16\].FF REGF\[25\].RFW.CG\[2\]/GCLK DW[16] VGND VGND VPWR VPWR
+ REGF\[25\].RFW.BIT\[16\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_48_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC1.D1.AND4 DEC1.D1.AND7/A DEC1.D1.AND7/B DEC1.D1.AND7/C DEC1.D1.AND7/D VGND VGND
+ VPWR VPWR DEC1.D1.AND4/X sky130_fd_sc_hd__and4bb_2
XREGF\[25\].RFW.BIT\[27\].OBUF2 REGF\[25\].RFW.BIT\[27\].FF/Q REGF\[25\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[27] sky130_fd_sc_hd__ebufn_2
Xfill_3_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[24\].RFW.CG\[3\] CLK REGF\[24\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[24\].RFW.CG\[3\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[26\].RFW.BIT\[6\].OBUF2 REGF\[26\].RFW.BIT\[6\].FF/Q REGF\[26\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[6] sky130_fd_sc_hd__ebufn_2
XREGF\[30\].RFW.BIT\[16\].OBUF2 REGF\[30\].RFW.BIT\[16\].FF/Q REGF\[30\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[16] sky130_fd_sc_hd__ebufn_2
Xfill_23_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_23_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[21\].RFW.BIT\[0\].OBUF1 REGF\[21\].RFW.BIT\[0\].FF/Q REGF\[21\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[0] sky130_fd_sc_hd__ebufn_2
Xtap_6_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.BIT\[3\].FF REGF\[18\].RFW.CG\[0\]/GCLK DW[3] VGND VGND VPWR VPWR
+ REGF\[18\].RFW.BIT\[3\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[2\].RFW.BIT\[19\].OBUF1 REGF\[2\].RFW.BIT\[19\].FF/Q REGF\[2\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[19] sky130_fd_sc_hd__ebufn_2
XREGF\[14\].RFW.BIT\[29\].FF REGF\[14\].RFW.CG\[3\]/GCLK DW[29] VGND VGND VPWR VPWR
+ REGF\[14\].RFW.BIT\[29\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[15\].RFW.BIT\[25\].OBUF1 REGF\[15\].RFW.BIT\[25\].FF/Q REGF\[15\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[25] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.BIT\[12\].OBUF2 REGF\[28\].RFW.BIT\[12\].FF/Q REGF\[28\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[12] sky130_fd_sc_hd__ebufn_2
XREGF\[10\].RFW.BIT\[31\].FF REGF\[10\].RFW.CG\[3\]/GCLK DW[31] VGND VGND VPWR VPWR
+ REGF\[10\].RFW.BIT\[31\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_20_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[14\].OBUF1 REGF\[20\].RFW.BIT\[14\].FF/Q REGF\[20\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[14] sky130_fd_sc_hd__ebufn_2
Xfill_48_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_48_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_48_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_6_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[17\].RFW.BIT\[5\].FF REGF\[17\].RFW.CG\[0\]/GCLK DW[5] VGND VGND VPWR VPWR
+ REGF\[17\].RFW.BIT\[5\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[18\].RFW.BIT\[10\].OBUF1 REGF\[18\].RFW.BIT\[10\].FF/Q REGF\[18\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[10] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.INV1\[2\] DEC0.D3.AND0/Y VGND VGND VPWR VPWR REGF\[24\].RFW.INV1\[2\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_13_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[23\].RFW.CG\[0\] CLK REGF\[23\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[23\].RFW.CG\[0\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XDEC0.D2.AND6 DEC0.D2.AND7/A DEC0.D2.AND7/B DEC0.D2.AND7/C DEC0.D2.AND7/D VGND VGND
+ VPWR VPWR DEC0.D2.AND6/X sky130_fd_sc_hd__and4b_2
XREGF\[19\].RFW.BIT\[26\].OBUF2 REGF\[19\].RFW.BIT\[26\].FF/Q REGF\[19\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[26] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[7\].FF REGF\[16\].RFW.CG\[0\]/GCLK DW[7] VGND VGND VPWR VPWR
+ REGF\[16\].RFW.BIT\[7\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_41_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[28\].RFW.BIT\[6\].OBUF2 REGF\[28\].RFW.BIT\[6\].FF/Q REGF\[28\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[6] sky130_fd_sc_hd__ebufn_2
XREGF\[11\].RFW.BIT\[28\].OBUF1 REGF\[11\].RFW.BIT\[28\].FF/Q REGF\[11\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[28] sky130_fd_sc_hd__ebufn_2
XREGF\[23\].RFW.BIT\[0\].OBUF1 REGF\[23\].RFW.BIT\[0\].FF/Q REGF\[23\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[0] sky130_fd_sc_hd__ebufn_2
Xfill_34_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[24\].RFW.BIT\[15\].OBUF2 REGF\[24\].RFW.BIT\[15\].FF/Q REGF\[24\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[15] sky130_fd_sc_hd__ebufn_2
Xfill_27_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_1_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XREGF\[30\].RFW.BIT\[9\].OBUF1 REGF\[30\].RFW.BIT\[9\].FF/Q REGF\[30\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[9] sky130_fd_sc_hd__ebufn_2
XREGF\[2\].RFW.BIT\[20\].OBUF1 REGF\[2\].RFW.BIT\[20\].FF/Q REGF\[2\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[20] sky130_fd_sc_hd__ebufn_2
XREGF\[14\].RFW.BIT\[13\].OBUF1 REGF\[14\].RFW.BIT\[13\].FF/Q REGF\[14\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[13] sky130_fd_sc_hd__ebufn_2
XREGF\[15\].RFW.BIT\[9\].FF REGF\[15\].RFW.CG\[1\]/GCLK DW[9] VGND VGND VPWR VPWR
+ REGF\[15\].RFW.BIT\[9\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[12\].RFW.CG\[3\] CLK REGF\[12\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[12\].RFW.CG\[3\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[21\].RFW.BIT\[4\].OBUF2 REGF\[21\].RFW.BIT\[4\].FF/Q REGF\[21\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[4] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[24\].FF REGF\[5\].RFW.CG\[3\]/GCLK DW[24] VGND VGND VPWR VPWR
+ REGF\[5\].RFW.BIT\[24\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[11\].RFW.BIT\[14\].FF REGF\[11\].RFW.CG\[1\]/GCLK DW[14] VGND VGND VPWR VPWR
+ REGF\[11\].RFW.BIT\[14\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_18_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[15\].RFW.BIT\[29\].OBUF2 REGF\[15\].RFW.BIT\[29\].FF/Q REGF\[15\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[29] sky130_fd_sc_hd__ebufn_2
Xfill_34_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[18\].OBUF2 REGF\[20\].RFW.BIT\[18\].FF/Q REGF\[20\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[18] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.BIT\[31\].OBUF2 REGF\[21\].RFW.BIT\[31\].FF/Q REGF\[21\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[31] sky130_fd_sc_hd__ebufn_2
Xfill_50_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_50_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_50_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[6\].RFW.BIT\[21\].OBUF2 REGF\[6\].RFW.BIT\[21\].FF/Q REGF\[6\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[21] sky130_fd_sc_hd__ebufn_2
XREGF\[25\].RFW.BIT\[0\].OBUF1 REGF\[25\].RFW.BIT\[0\].FF/Q REGF\[25\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[0] sky130_fd_sc_hd__ebufn_2
Xfill_59_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_59_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_59_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_59_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_59_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.BIT\[14\].OBUF2 REGF\[18\].RFW.BIT\[14\].FF/Q REGF\[18\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[14] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.BIT\[7\].FF REGF\[29\].RFW.CG\[0\]/GCLK DW[7] VGND VGND VPWR VPWR
+ REGF\[29\].RFW.BIT\[7\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_11_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[10\].RFW.BIT\[16\].OBUF1 REGF\[10\].RFW.BIT\[16\].FF/Q REGF\[10\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[16] sky130_fd_sc_hd__ebufn_2
XREGF\[22\].RFW.BIT\[24\].FF REGF\[22\].RFW.CG\[3\]/GCLK DW[24] VGND VGND VPWR VPWR
+ REGF\[22\].RFW.BIT\[24\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[11\].RFW.CG\[0\] CLK REGF\[11\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[11\].RFW.CG\[0\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[19\].RFW.INV1\[3\] DEC0.D2.AND3/X VGND VGND VPWR VPWR REGF\[19\].RFW.INV1\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[23\].RFW.BIT\[4\].OBUF2 REGF\[23\].RFW.BIT\[4\].FF/Q REGF\[23\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[4] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.BIT\[9\].FF REGF\[28\].RFW.CG\[1\]/GCLK DW[9] VGND VGND VPWR VPWR
+ REGF\[28\].RFW.BIT\[9\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[17\].RFW.BIT\[31\].FF REGF\[17\].RFW.CG\[3\]/GCLK DW[31] VGND VGND VPWR VPWR
+ REGF\[17\].RFW.BIT\[31\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[2\].RFW.BIT\[24\].OBUF2 REGF\[2\].RFW.BIT\[24\].FF/Q REGF\[2\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[24] sky130_fd_sc_hd__ebufn_2
Xfill_32_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[14\].RFW.BIT\[17\].OBUF2 REGF\[14\].RFW.BIT\[17\].FF/Q REGF\[14\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[17] sky130_fd_sc_hd__ebufn_2
XREGF\[15\].RFW.BIT\[30\].OBUF2 REGF\[15\].RFW.BIT\[30\].FF/Q REGF\[15\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[30] sky130_fd_sc_hd__ebufn_2
Xfill_25_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_18_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XDEC1.D0.ABUF\[2\] RB[2] VGND VGND VPWR VPWR DEC1.D0.AND7/C sky130_fd_sc_hd__clkbuf_2
XREGF\[27\].RFW.BIT\[0\].OBUF1 REGF\[27\].RFW.BIT\[0\].FF/Q REGF\[27\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[0] sky130_fd_sc_hd__ebufn_2
Xfill_20_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_29_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_29_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_29_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_45_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_45_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_45_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[25\].RFW.BIT\[4\].OBUF2 REGF\[25\].RFW.BIT\[4\].FF/Q REGF\[25\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[4] sky130_fd_sc_hd__ebufn_2
Xfill_45_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_61_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_61_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_61_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_61_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_61_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_59_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_10_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[1\].RFW.BIT\[12\].OBUF2 REGF\[1\].RFW.BIT\[12\].FF/Q REGF\[1\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[12] sky130_fd_sc_hd__ebufn_2
Xfill_19_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.BIT\[14\].FF REGF\[18\].RFW.CG\[1\]/GCLK DW[14] VGND VGND VPWR VPWR
+ REGF\[18\].RFW.BIT\[14\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_19_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[29\].RFW.BIT\[0\].OBUF1 REGF\[29\].RFW.BIT\[0\].FF/Q REGF\[29\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[0] sky130_fd_sc_hd__ebufn_2
Xfill_11_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_35_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.BIT\[19\].OBUF1 REGF\[31\].RFW.BIT\[19\].FF/Q REGF\[31\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[19] sky130_fd_sc_hd__ebufn_2
Xfill_7_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_7_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_7_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[29\].RFW.BIT\[15\].OBUF1 REGF\[29\].RFW.BIT\[15\].FF/Q REGF\[29\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[15] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[4\].OBUF2 REGF\[27\].RFW.BIT\[4\].FF/Q REGF\[27\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[4] sky130_fd_sc_hd__ebufn_2
Xfill_30_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[29\].RFW.BIT\[24\].FF REGF\[29\].RFW.CG\[3\]/GCLK DW[24] VGND VGND VPWR VPWR
+ REGF\[29\].RFW.BIT\[24\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[6\].RFW.INV1\[1\] DEC0.D0.AND6/X VGND VGND VPWR VPWR REGF\[6\].RFW.INV1\[1\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_15_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[10\].RFW.BIT\[21\].OBUF2 REGF\[10\].RFW.BIT\[21\].FF/Q REGF\[10\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[21] sky130_fd_sc_hd__ebufn_2
Xfill_31_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_52_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_31_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[2\].OBUF2 REGF\[20\].RFW.BIT\[2\].FF/Q REGF\[20\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[2] sky130_fd_sc_hd__ebufn_2
Xtap_38_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_56_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_56_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_56_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[25\].RFW.BIT\[18\].OBUF1 REGF\[25\].RFW.BIT\[18\].FF/Q REGF\[25\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[18] sky130_fd_sc_hd__ebufn_2
XREGF\[3\].RFW.BIT\[15\].FF REGF\[3\].RFW.CG\[1\]/GCLK DW[15] VGND VGND VPWR VPWR
+ REGF\[3\].RFW.BIT\[15\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[26\].RFW.BIT\[31\].OBUF1 REGF\[26\].RFW.BIT\[31\].FF/Q REGF\[26\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[31] sky130_fd_sc_hd__ebufn_2
XDEC2.D3.AND0 DEC2.D3.AND7/A DEC2.D3.AND7/B DEC2.D3.AND7/C DEC2.D3.AND7/D VGND VGND
+ VPWR VPWR DEC2.D3.AND0/Y sky130_fd_sc_hd__nor4b_2
XREGF\[31\].RFW.BIT\[20\].OBUF1 REGF\[31\].RFW.BIT\[20\].FF/Q REGF\[31\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[20] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.BIT\[4\].OBUF2 REGF\[29\].RFW.BIT\[4\].FF/Q REGF\[29\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[4] sky130_fd_sc_hd__ebufn_2
Xfill_21_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_21_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfill_59_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.BIT\[7\].OBUF1 REGF\[31\].RFW.BIT\[7\].FF/Q REGF\[31\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[7] sky130_fd_sc_hd__ebufn_2
XREGF\[20\].RFW.BIT\[15\].FF REGF\[20\].RFW.CG\[1\]/GCLK DW[15] VGND VGND VPWR VPWR
+ REGF\[20\].RFW.BIT\[15\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_7_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[29\].RFW.BIT\[19\].OBUF2 REGF\[29\].RFW.BIT\[19\].FF/Q REGF\[29\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[19] sky130_fd_sc_hd__ebufn_2
XREGF\[22\].RFW.BIT\[2\].OBUF2 REGF\[22\].RFW.BIT\[2\].FF/Q REGF\[22\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[2] sky130_fd_sc_hd__ebufn_2
XREGF\[13\].RFW.BIT\[0\].FF REGF\[13\].RFW.CG\[0\]/GCLK DW[0] VGND VGND VPWR VPWR
+ REGF\[13\].RFW.BIT\[0\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[7\].RFW.BIT\[24\].OBUF1 REGF\[7\].RFW.BIT\[24\].FF/Q REGF\[7\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[24] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.BIT\[17\].OBUF1 REGF\[19\].RFW.BIT\[17\].FF/Q REGF\[19\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[17] sky130_fd_sc_hd__ebufn_2
Xtap_0_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[15\].RFW.BIT\[22\].FF REGF\[15\].RFW.CG\[2\]/GCLK DW[22] VGND VGND VPWR VPWR
+ REGF\[15\].RFW.BIT\[22\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_26_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[12\].RFW.BIT\[2\].FF REGF\[12\].RFW.CG\[0\]/GCLK DW[2] VGND VGND VPWR VPWR
+ REGF\[12\].RFW.BIT\[2\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[31\].RFW.BIT\[25\].FF REGF\[31\].RFW.CG\[3\]/GCLK DW[25] VGND VGND VPWR VPWR
+ REGF\[31\].RFW.BIT\[25\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_42_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_42_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_42_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_50_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_43_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_36_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[11\].RFW.BIT\[4\].FF REGF\[11\].RFW.CG\[0\]/GCLK DW[4] VGND VGND VPWR VPWR
+ REGF\[11\].RFW.BIT\[4\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[31\].RFW.BIT\[24\].OBUF2 REGF\[31\].RFW.BIT\[24\].FF/Q REGF\[31\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[24] sky130_fd_sc_hd__ebufn_2
XREGF\[20\].RFW.INV2\[0\] DEC1.D2.AND4/X VGND VGND VPWR VPWR REGF\[20\].RFW.INV2\[0\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[24\].RFW.BIT\[2\].OBUF2 REGF\[24\].RFW.BIT\[2\].FF/Q REGF\[24\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[2] sky130_fd_sc_hd__ebufn_2
XREGF\[3\].RFW.BIT\[27\].OBUF1 REGF\[3\].RFW.BIT\[27\].FF/Q REGF\[3\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[27] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.BIT\[20\].OBUF2 REGF\[29\].RFW.BIT\[20\].FF/Q REGF\[29\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[20] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.BIT\[22\].OBUF1 REGF\[21\].RFW.BIT\[22\].FF/Q REGF\[21\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[22] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[0\].FF REGF\[26\].RFW.CG\[0\]/GCLK DW[0] VGND VGND VPWR VPWR
+ REGF\[26\].RFW.BIT\[0\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[10\].RFW.BIT\[6\].FF REGF\[10\].RFW.CG\[0\]/GCLK DW[6] VGND VGND VPWR VPWR
+ REGF\[10\].RFW.BIT\[6\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[6\].RFW.BIT\[12\].OBUF1 REGF\[6\].RFW.BIT\[12\].FF/Q REGF\[6\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[12] sky130_fd_sc_hd__ebufn_2
Xfill_57_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_4_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_4_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[25\].RFW.BIT\[2\].FF REGF\[25\].RFW.CG\[0\]/GCLK DW[2] VGND VGND VPWR VPWR
+ REGF\[25\].RFW.BIT\[2\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[9\].RFW.CG\[2\] CLK REGF\[9\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[9\].RFW.CG\[2\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[20\].RFW.CG\[2\] CLK REGF\[20\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[20\].RFW.CG\[2\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_5_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[7\].RFW.BIT\[28\].OBUF2 REGF\[7\].RFW.BIT\[28\].FF/Q REGF\[7\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[28] sky130_fd_sc_hd__ebufn_2
XREGF\[25\].RFW.BIT\[23\].OBUF2 REGF\[25\].RFW.BIT\[23\].FF/Q REGF\[25\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[23] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[4\].FF REGF\[24\].RFW.CG\[0\]/GCLK DW[4] VGND VGND VPWR VPWR
+ REGF\[24\].RFW.BIT\[4\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[30\].RFW.BIT\[12\].OBUF2 REGF\[30\].RFW.BIT\[12\].FF/Q REGF\[30\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[12] sky130_fd_sc_hd__ebufn_2
Xtap_22_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[26\].RFW.BIT\[2\].OBUF2 REGF\[26\].RFW.BIT\[2\].FF/Q REGF\[26\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[2] sky130_fd_sc_hd__ebufn_2
XREGF\[2\].RFW.BIT\[15\].OBUF1 REGF\[2\].RFW.BIT\[15\].FF/Q REGF\[2\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[15] sky130_fd_sc_hd__ebufn_2
Xfill_37_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_37_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_37_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xtap_8_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[15\].RFW.BIT\[21\].OBUF1 REGF\[15\].RFW.BIT\[21\].FF/Q REGF\[15\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[21] sky130_fd_sc_hd__ebufn_2
Xtap_14_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_53_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_53_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_53_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_53_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[27\].RFW.BIT\[15\].FF REGF\[27\].RFW.CG\[1\]/GCLK DW[15] VGND VGND VPWR VPWR
+ REGF\[27\].RFW.BIT\[15\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[20\].RFW.BIT\[10\].OBUF1 REGF\[20\].RFW.BIT\[10\].FF/Q REGF\[20\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[10] sky130_fd_sc_hd__ebufn_2
XDEC2.D0.AND3 DEC2.D0.AND7/C DEC2.D0.AND7/B DEC2.D0.AND7/A DEC2.D0.AND7/D VGND VGND
+ VPWR VPWR DEC2.D0.AND3/X sky130_fd_sc_hd__and4b_2
XREGF\[23\].RFW.BIT\[6\].FF REGF\[23\].RFW.CG\[0\]/GCLK DW[6] VGND VGND VPWR VPWR
+ REGF\[23\].RFW.BIT\[6\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_41_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[15\].RFW.INV2\[1\] DEC1.D1.AND7/X VGND VGND VPWR VPWR REGF\[15\].RFW.INV2\[1\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[21\].RFW.BIT\[26\].OBUF2 REGF\[21\].RFW.BIT\[26\].FF/Q REGF\[21\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[26] sky130_fd_sc_hd__ebufn_2
XREGF\[9\].RFW.BIT\[1\].FF REGF\[9\].RFW.CG\[0\]/GCLK DW[1] VGND VGND VPWR VPWR REGF\[9\].RFW.BIT\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[16\].RFW.BIT\[28\].FF REGF\[16\].RFW.CG\[3\]/GCLK DW[28] VGND VGND VPWR VPWR
+ REGF\[16\].RFW.BIT\[28\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[12\].RFW.BIT\[30\].FF REGF\[12\].RFW.CG\[3\]/GCLK DW[30] VGND VGND VPWR VPWR
+ REGF\[12\].RFW.BIT\[30\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_27_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_27_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_29_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[22\].RFW.BIT\[8\].FF REGF\[22\].RFW.CG\[1\]/GCLK DW[8] VGND VGND VPWR VPWR
+ REGF\[22\].RFW.BIT\[8\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[6\].RFW.BIT\[16\].OBUF2 REGF\[6\].RFW.BIT\[16\].FF/Q REGF\[6\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[16] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.BIT\[22\].OBUF2 REGF\[19\].RFW.BIT\[22\].FF/Q REGF\[19\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[22] sky130_fd_sc_hd__ebufn_2
Xfill_43_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[28\].RFW.BIT\[2\].OBUF2 REGF\[28\].RFW.BIT\[2\].FF/Q REGF\[28\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[2] sky130_fd_sc_hd__ebufn_2
XREGF\[11\].RFW.BIT\[24\].OBUF1 REGF\[11\].RFW.BIT\[24\].FF/Q REGF\[11\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[24] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[11\].OBUF2 REGF\[24\].RFW.BIT\[11\].FF/Q REGF\[24\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[11] sky130_fd_sc_hd__ebufn_2
XREGF\[8\].RFW.BIT\[3\].FF REGF\[8\].RFW.CG\[0\]/GCLK DW[3] VGND VGND VPWR VPWR REGF\[8\].RFW.BIT\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xfill_62_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_55_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[30\].RFW.BIT\[5\].OBUF1 REGF\[30\].RFW.BIT\[5\].FF/Q REGF\[30\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[5] sky130_fd_sc_hd__ebufn_2
XDEC1.D1.AND5 DEC1.D1.AND7/B DEC1.D1.AND7/A DEC1.D1.AND7/C DEC1.D1.AND7/D VGND VGND
+ VPWR VPWR DEC1.D1.AND5/X sky130_fd_sc_hd__and4b_2
Xfill_48_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDEC2.D3.ABUF\[1\] RW[1] VGND VGND VPWR VPWR DEC2.D3.AND7/B sky130_fd_sc_hd__clkbuf_2
Xfill_3_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[7\].RFW.BIT\[5\].FF REGF\[7\].RFW.CG\[0\]/GCLK DW[5] VGND VGND VPWR VPWR REGF\[7\].RFW.BIT\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xfill_23_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[21\].RFW.BIT\[0\].OBUF2 REGF\[21\].RFW.BIT\[0\].FF/Q REGF\[21\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[0] sky130_fd_sc_hd__ebufn_2
XREGF\[11\].RFW.INV1\[2\] DEC0.D1.AND3/X VGND VGND VPWR VPWR REGF\[11\].RFW.INV1\[2\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[2\].RFW.BIT\[19\].OBUF2 REGF\[2\].RFW.BIT\[19\].FF/Q REGF\[2\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[19] sky130_fd_sc_hd__ebufn_2
XREGF\[15\].RFW.BIT\[25\].OBUF2 REGF\[15\].RFW.BIT\[25\].FF/Q REGF\[15\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[25] sky130_fd_sc_hd__ebufn_2
Xtap_20_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[27\].RFW.INV1\[3\] DEC0.D3.AND3/X VGND VGND VPWR VPWR REGF\[27\].RFW.INV1\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[20\].RFW.BIT\[14\].OBUF2 REGF\[20\].RFW.BIT\[14\].FF/Q REGF\[20\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[14] sky130_fd_sc_hd__ebufn_2
Xfill_48_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_48_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_48_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[6\].RFW.BIT\[7\].FF REGF\[6\].RFW.CG\[0\]/GCLK DW[7] VGND VGND VPWR VPWR REGF\[6\].RFW.BIT\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xtap_6_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[1\].RFW.BIT\[29\].FF REGF\[1\].RFW.CG\[3\]/GCLK DW[29] VGND VGND VPWR VPWR
+ REGF\[1\].RFW.BIT\[29\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[7\].RFW.BIT\[23\].FF REGF\[7\].RFW.CG\[2\]/GCLK DW[23] VGND VGND VPWR VPWR
+ REGF\[7\].RFW.BIT\[23\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[13\].RFW.BIT\[13\].FF REGF\[13\].RFW.CG\[1\]/GCLK DW[13] VGND VGND VPWR VPWR
+ REGF\[13\].RFW.BIT\[13\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[18\].RFW.BIT\[10\].OBUF2 REGF\[18\].RFW.BIT\[10\].FF/Q REGF\[18\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[10] sky130_fd_sc_hd__ebufn_2
XREGF\[10\].RFW.BIT\[12\].OBUF1 REGF\[10\].RFW.BIT\[12\].FF/Q REGF\[10\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[12] sky130_fd_sc_hd__ebufn_2
Xfill_13_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_13_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_13_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_13_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC0.D2.AND7 DEC0.D2.AND7/A DEC0.D2.AND7/B DEC0.D2.AND7/C DEC0.D2.AND7/D VGND VGND
+ VPWR VPWR DEC0.D2.AND7/X sky130_fd_sc_hd__and4_2
XREGF\[5\].RFW.BIT\[9\].FF REGF\[5\].RFW.CG\[1\]/GCLK DW[9] VGND VGND VPWR VPWR REGF\[5\].RFW.BIT\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xfill_41_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[11\].RFW.BIT\[28\].OBUF2 REGF\[11\].RFW.BIT\[28\].FF/Q REGF\[11\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[28] sky130_fd_sc_hd__ebufn_2
XREGF\[23\].RFW.BIT\[0\].OBUF2 REGF\[23\].RFW.BIT\[0\].FF/Q REGF\[23\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[0] sky130_fd_sc_hd__ebufn_2
Xfill_34_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_27_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_1_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_1_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_1_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[24\].RFW.BIT\[23\].FF REGF\[24\].RFW.CG\[2\]/GCLK DW[23] VGND VGND VPWR VPWR
+ REGF\[24\].RFW.BIT\[23\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[30\].RFW.BIT\[9\].OBUF2 REGF\[30\].RFW.BIT\[9\].FF/Q REGF\[30\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[9] sky130_fd_sc_hd__ebufn_2
XREGF\[2\].RFW.BIT\[20\].OBUF2 REGF\[2\].RFW.BIT\[20\].FF/Q REGF\[2\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[20] sky130_fd_sc_hd__ebufn_2
XREGF\[14\].RFW.BIT\[13\].OBUF2 REGF\[14\].RFW.BIT\[13\].FF/Q REGF\[14\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[13] sky130_fd_sc_hd__ebufn_2
Xfill_60_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_18_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[19\].RFW.BIT\[30\].FF REGF\[19\].RFW.CG\[3\]/GCLK DW[30] VGND VGND VPWR VPWR
+ REGF\[19\].RFW.BIT\[30\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_50_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_50_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_50_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[25\].RFW.BIT\[0\].OBUF2 REGF\[25\].RFW.BIT\[0\].FF/Q REGF\[25\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[0] sky130_fd_sc_hd__ebufn_2
Xfill_59_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_59_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_59_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_59_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_11_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[10\].RFW.BIT\[16\].OBUF2 REGF\[10\].RFW.BIT\[16\].FF/Q REGF\[10\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[16] sky130_fd_sc_hd__ebufn_2
Xtap_4_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[26\].RFW.BIT\[26\].OBUF1 REGF\[26\].RFW.BIT\[26\].FF/Q REGF\[26\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[26] sky130_fd_sc_hd__ebufn_2
XREGF\[31\].RFW.BIT\[15\].OBUF1 REGF\[31\].RFW.BIT\[15\].FF/Q REGF\[31\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[15] sky130_fd_sc_hd__ebufn_2
Xfill_32_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_25_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[8\].RFW.BIT\[29\].FF REGF\[8\].RFW.CG\[3\]/GCLK DW[29] VGND VGND VPWR VPWR
+ REGF\[8\].RFW.BIT\[29\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[14\].RFW.BIT\[19\].FF REGF\[14\].RFW.CG\[2\]/GCLK DW[19] VGND VGND VPWR VPWR
+ REGF\[14\].RFW.BIT\[19\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_18_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XREGF\[29\].RFW.BIT\[11\].OBUF1 REGF\[29\].RFW.BIT\[11\].FF/Q REGF\[29\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[11] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.BIT\[31\].FF REGF\[4\].RFW.CG\[3\]/GCLK DW[31] VGND VGND VPWR VPWR
+ REGF\[4\].RFW.BIT\[31\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[10\].RFW.BIT\[21\].FF REGF\[10\].RFW.CG\[2\]/GCLK DW[21] VGND VGND VPWR VPWR
+ REGF\[10\].RFW.BIT\[21\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[27\].RFW.BIT\[0\].OBUF2 REGF\[27\].RFW.BIT\[0\].FF/Q REGF\[27\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[0] sky130_fd_sc_hd__ebufn_2
Xfill_29_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_29_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[22\].RFW.BIT\[29\].OBUF1 REGF\[22\].RFW.BIT\[29\].FF/Q REGF\[22\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[29] sky130_fd_sc_hd__ebufn_2
Xfill_45_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_45_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_45_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XREGF\[7\].RFW.BIT\[19\].OBUF1 REGF\[7\].RFW.BIT\[19\].FF/Q REGF\[7\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[19] sky130_fd_sc_hd__ebufn_2
Xtap_22_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[25\].RFW.BIT\[29\].FF REGF\[25\].RFW.CG\[3\]/GCLK DW[29] VGND VGND VPWR VPWR
+ REGF\[25\].RFW.BIT\[29\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_61_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_61_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_61_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_61_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[21\].RFW.BIT\[31\].FF REGF\[21\].RFW.CG\[3\]/GCLK DW[31] VGND VGND VPWR VPWR
+ REGF\[21\].RFW.BIT\[31\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_59_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[25\].RFW.BIT\[14\].OBUF1 REGF\[25\].RFW.BIT\[14\].FF/Q REGF\[25\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[14] sky130_fd_sc_hd__ebufn_2
Xfill_10_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_10_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_19_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_19_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[29\].RFW.BIT\[0\].OBUF2 REGF\[29\].RFW.BIT\[0\].FF/Q REGF\[29\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[0] sky130_fd_sc_hd__ebufn_2
Xfill_11_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.BIT\[19\].OBUF2 REGF\[31\].RFW.BIT\[19\].FF/Q REGF\[31\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[19] sky130_fd_sc_hd__ebufn_2
XREGF\[31\].RFW.BIT\[3\].OBUF1 REGF\[31\].RFW.BIT\[3\].FF/Q REGF\[31\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[3] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[14\].FF REGF\[5\].RFW.CG\[1\]/GCLK DW[14] VGND VGND VPWR VPWR
+ REGF\[5\].RFW.BIT\[14\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_51_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[9\].RFW.INV1\[2\] DEC0.D1.AND1/X VGND VGND VPWR VPWR REGF\[9\].RFW.INV1\[2\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_7_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_7_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_7_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_7_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[16\].RFW.BIT\[28\].OBUF1 REGF\[16\].RFW.BIT\[28\].FF/Q REGF\[16\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[28] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.BIT\[15\].OBUF2 REGF\[29\].RFW.BIT\[15\].FF/Q REGF\[29\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[15] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.BIT\[17\].OBUF1 REGF\[21\].RFW.BIT\[17\].FF/Q REGF\[21\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[17] sky130_fd_sc_hd__ebufn_2
XREGF\[22\].RFW.BIT\[30\].OBUF1 REGF\[22\].RFW.BIT\[30\].FF/Q REGF\[22\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[30] sky130_fd_sc_hd__ebufn_2
Xfill_30_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_23_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[7\].RFW.BIT\[20\].OBUF1 REGF\[7\].RFW.BIT\[20\].FF/Q REGF\[7\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[20] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.BIT\[13\].OBUF1 REGF\[19\].RFW.BIT\[13\].FF/Q REGF\[19\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[13] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.INV1\[0\] DEC0.D3.AND5/X VGND VGND VPWR VPWR REGF\[29\].RFW.INV1\[0\]/Y
+ sky130_fd_sc_hd__inv_4
Xtap_52_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[22\].RFW.BIT\[14\].FF REGF\[22\].RFW.CG\[1\]/GCLK DW[14] VGND VGND VPWR VPWR
+ REGF\[22\].RFW.BIT\[14\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_31_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_38_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_56_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_56_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_56_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[25\].RFW.BIT\[18\].OBUF2 REGF\[25\].RFW.BIT\[18\].FF/Q REGF\[25\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[18] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[31\].OBUF2 REGF\[26\].RFW.BIT\[31\].FF/Q REGF\[26\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[31] sky130_fd_sc_hd__ebufn_2
XREGF\[11\].RFW.BIT\[27\].FF REGF\[11\].RFW.CG\[3\]/GCLK DW[27] VGND VGND VPWR VPWR
+ REGF\[11\].RFW.BIT\[27\].FF/Q sky130_fd_sc_hd__dfxtp_1
XDEC2.D3.AND1 DEC2.D3.AND7/C DEC2.D3.AND7/B DEC2.D3.AND7/A DEC2.D3.AND7/D VGND VGND
+ VPWR VPWR DEC2.D3.AND1/X sky130_fd_sc_hd__and4bb_2
XREGF\[31\].RFW.BIT\[20\].OBUF2 REGF\[31\].RFW.BIT\[20\].FF/Q REGF\[31\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[20] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.BIT\[21\].FF REGF\[17\].RFW.CG\[2\]/GCLK DW[21] VGND VGND VPWR VPWR
+ REGF\[17\].RFW.BIT\[21\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_21_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.BIT\[0\].FF REGF\[3\].RFW.CG\[0\]/GCLK DW[0] VGND VGND VPWR VPWR REGF\[3\].RFW.BIT\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[3\].RFW.BIT\[23\].OBUF1 REGF\[3\].RFW.BIT\[23\].FF/Q REGF\[3\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[23] sky130_fd_sc_hd__ebufn_2
Xfill_21_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[15\].RFW.BIT\[16\].OBUF1 REGF\[15\].RFW.BIT\[16\].FF/Q REGF\[15\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[16] sky130_fd_sc_hd__ebufn_2
Xfill_59_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[31\].RFW.BIT\[7\].OBUF2 REGF\[31\].RFW.BIT\[7\].FF/Q REGF\[31\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[7] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.CG\[1\] CLK REGF\[5\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[5\].RFW.CG\[1\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_7_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[31\].RFW.BIT\[3\].FF REGF\[31\].RFW.CG\[0\]/GCLK DW[3] VGND VGND VPWR VPWR
+ REGF\[31\].RFW.BIT\[3\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[2\].RFW.BIT\[2\].FF REGF\[2\].RFW.CG\[0\]/GCLK DW[2] VGND VGND VPWR VPWR REGF\[2\].RFW.BIT\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[28\].RFW.BIT\[31\].FF REGF\[28\].RFW.CG\[3\]/GCLK DW[31] VGND VGND VPWR VPWR
+ REGF\[28\].RFW.BIT\[31\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[31\].RFW.CGAND DEC2.D3.AND7/X WE VGND VGND VPWR VPWR REGF\[31\].RFW.CGAND/X
+ sky130_fd_sc_hd__and2_1
XREGF\[3\].RFW.INV2\[3\] DEC1.D0.AND3/X VGND VGND VPWR VPWR REGF\[3\].RFW.INV2\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[7\].RFW.BIT\[24\].OBUF2 REGF\[7\].RFW.BIT\[24\].FF/Q REGF\[7\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[24] sky130_fd_sc_hd__ebufn_2
Xtap_0_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[19\].RFW.BIT\[17\].OBUF2 REGF\[19\].RFW.BIT\[17\].FF/Q REGF\[19\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[17] sky130_fd_sc_hd__ebufn_2
XREGF\[30\].RFW.BIT\[5\].FF REGF\[30\].RFW.CG\[0\]/GCLK DW[5] VGND VGND VPWR VPWR
+ REGF\[30\].RFW.BIT\[5\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[1\].RFW.BIT\[4\].FF REGF\[1\].RFW.CG\[0\]/GCLK DW[4] VGND VGND VPWR VPWR REGF\[1\].RFW.BIT\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[11\].RFW.BIT\[19\].OBUF1 REGF\[11\].RFW.BIT\[19\].FF/Q REGF\[11\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[19] sky130_fd_sc_hd__ebufn_2
Xfill_26_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_42_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[2\].RFW.BIT\[22\].FF REGF\[2\].RFW.CG\[2\]/GCLK DW[22] VGND VGND VPWR VPWR
+ REGF\[2\].RFW.BIT\[22\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[2\].RFW.BIT\[11\].OBUF1 REGF\[2\].RFW.BIT\[11\].FF/Q REGF\[2\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[11] sky130_fd_sc_hd__ebufn_2
XREGF\[23\].RFW.INV2\[1\] DEC1.D2.AND7/X VGND VGND VPWR VPWR REGF\[23\].RFW.INV2\[1\]/Y
+ sky130_fd_sc_hd__inv_4
Xtap_50_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_36_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.BIT\[27\].OBUF2 REGF\[3\].RFW.BIT\[27\].FF/Q REGF\[3\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[27] sky130_fd_sc_hd__ebufn_2
Xfill_16_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[21\].RFW.BIT\[22\].OBUF2 REGF\[21\].RFW.BIT\[22\].FF/Q REGF\[21\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[22] sky130_fd_sc_hd__ebufn_2
Xfill_32_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[6\].RFW.BIT\[12\].OBUF2 REGF\[6\].RFW.BIT\[12\].FF/Q REGF\[6\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[12] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.BIT\[14\].FF REGF\[29\].RFW.CG\[1\]/GCLK DW[14] VGND VGND VPWR VPWR
+ REGF\[29\].RFW.BIT\[14\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_57_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_4_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_4_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_4_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[11\].RFW.BIT\[20\].OBUF1 REGF\[11\].RFW.BIT\[20\].FF/Q REGF\[11\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[20] sky130_fd_sc_hd__ebufn_2
Xfill_5_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[19\].RFW.CG\[0\] CLK REGF\[19\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[19\].RFW.CG\[0\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[30\].RFW.BIT\[1\].OBUF1 REGF\[30\].RFW.BIT\[1\].FF/Q REGF\[30\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[1] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.BIT\[27\].FF REGF\[18\].RFW.CG\[3\]/GCLK DW[27] VGND VGND VPWR VPWR
+ REGF\[18\].RFW.BIT\[27\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_22_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[2\].RFW.BIT\[15\].OBUF2 REGF\[2\].RFW.BIT\[15\].FF/Q REGF\[2\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[15] sky130_fd_sc_hd__ebufn_2
Xfill_37_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_37_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xtap_8_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_53_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_53_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[15\].RFW.BIT\[21\].OBUF2 REGF\[15\].RFW.BIT\[21\].FF/Q REGF\[15\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[21] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.INV2\[2\] DEC1.D2.AND2/X VGND VGND VPWR VPWR REGF\[18\].RFW.INV2\[2\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_53_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XREGF\[20\].RFW.BIT\[10\].OBUF2 REGF\[20\].RFW.BIT\[10\].FF/Q REGF\[20\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[10] sky130_fd_sc_hd__ebufn_2
XDEC2.D0.AND4 DEC2.D0.AND7/A DEC2.D0.AND7/B DEC2.D0.AND7/C DEC2.D0.AND7/D VGND VGND
+ VPWR VPWR DEC2.D0.AND4/X sky130_fd_sc_hd__and4bb_2
Xtap_30_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_41_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_27_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_27_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_43_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_43_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.BIT\[28\].FF REGF\[3\].RFW.CG\[3\]/GCLK DW[28] VGND VGND VPWR VPWR
+ REGF\[3\].RFW.BIT\[28\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[11\].RFW.BIT\[24\].OBUF2 REGF\[11\].RFW.BIT\[24\].FF/Q REGF\[11\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[24] sky130_fd_sc_hd__ebufn_2
XREGF\[9\].RFW.BIT\[22\].FF REGF\[9\].RFW.CG\[2\]/GCLK DW[22] VGND VGND VPWR VPWR
+ REGF\[9\].RFW.BIT\[22\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[15\].RFW.BIT\[12\].FF REGF\[15\].RFW.CG\[1\]/GCLK DW[12] VGND VGND VPWR VPWR
+ REGF\[15\].RFW.BIT\[12\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[31\].RFW.BIT\[15\].FF REGF\[31\].RFW.CG\[1\]/GCLK DW[15] VGND VGND VPWR VPWR
+ REGF\[31\].RFW.BIT\[15\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_62_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[30\].RFW.BIT\[5\].OBUF2 REGF\[30\].RFW.BIT\[5\].FF/Q REGF\[30\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[5] sky130_fd_sc_hd__ebufn_2
Xfill_55_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[14\].RFW.INV1\[3\] DEC0.D1.AND6/X VGND VGND VPWR VPWR REGF\[14\].RFW.INV1\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XDEC1.D1.AND6 DEC1.D1.AND7/A DEC1.D1.AND7/B DEC1.D1.AND7/C DEC1.D1.AND7/D VGND VGND
+ VPWR VPWR DEC1.D1.AND6/X sky130_fd_sc_hd__and4b_2
Xfill_48_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_3_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XREGF\[20\].RFW.BIT\[28\].FF REGF\[20\].RFW.CG\[3\]/GCLK DW[28] VGND VGND VPWR VPWR
+ REGF\[20\].RFW.BIT\[28\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[26\].RFW.BIT\[22\].FF REGF\[26\].RFW.CG\[2\]/GCLK DW[22] VGND VGND VPWR VPWR
+ REGF\[26\].RFW.BIT\[22\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_20_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_48_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_13_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_48_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_48_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[10\].RFW.BIT\[12\].OBUF2 REGF\[10\].RFW.BIT\[12\].FF/Q REGF\[10\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[12] sky130_fd_sc_hd__ebufn_2
Xfill_13_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_13_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_13_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC2.D1.ABUF\[0\] RW[0] VGND VGND VPWR VPWR DEC2.D1.AND7/A sky130_fd_sc_hd__clkbuf_2
Xfill_13_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XREGF\[8\].RFW.BIT\[27\].OBUF1 REGF\[8\].RFW.BIT\[27\].FF/Q REGF\[8\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[27] sky130_fd_sc_hd__ebufn_2
Xfill_41_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_34_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_27_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[26\].RFW.BIT\[22\].OBUF1 REGF\[26\].RFW.BIT\[22\].FF/Q REGF\[26\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[22] sky130_fd_sc_hd__ebufn_2
Xfill_1_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_1_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[31\].RFW.BIT\[11\].OBUF1 REGF\[31\].RFW.BIT\[11\].FF/Q REGF\[31\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[11] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.INV2\[0\] DEC1.D0.AND5/X VGND VGND VPWR VPWR REGF\[5\].RFW.INV2\[0\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_60_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_53_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[22\].RFW.BIT\[25\].OBUF1 REGF\[22\].RFW.BIT\[25\].FF/Q REGF\[22\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[25] sky130_fd_sc_hd__ebufn_2
Xfill_50_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[16\].RFW.BIT\[18\].FF REGF\[16\].RFW.CG\[2\]/GCLK DW[18] VGND VGND VPWR VPWR
+ REGF\[16\].RFW.BIT\[18\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_59_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.BIT\[30\].FF REGF\[6\].RFW.CG\[3\]/GCLK DW[30] VGND VGND VPWR VPWR
+ REGF\[6\].RFW.BIT\[30\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[12\].RFW.BIT\[20\].FF REGF\[12\].RFW.CG\[2\]/GCLK DW[20] VGND VGND VPWR VPWR
+ REGF\[12\].RFW.BIT\[20\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_59_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_59_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_59_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[7\].RFW.BIT\[15\].OBUF1 REGF\[7\].RFW.BIT\[15\].FF/Q REGF\[7\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[15] sky130_fd_sc_hd__ebufn_2
Xtap_11_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[25\].RFW.BIT\[10\].OBUF1 REGF\[25\].RFW.BIT\[10\].FF/Q REGF\[25\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[10] sky130_fd_sc_hd__ebufn_2
XREGF\[1\].RFW.INV1\[1\] DEC0.D0.AND1/X VGND VGND VPWR VPWR REGF\[1\].RFW.INV1\[1\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_24_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[26\].RFW.BIT\[26\].OBUF2 REGF\[26\].RFW.BIT\[26\].FF/Q REGF\[26\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[26] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[28\].FF REGF\[27\].RFW.CG\[3\]/GCLK DW[28] VGND VGND VPWR VPWR
+ REGF\[27\].RFW.BIT\[28\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_40_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[23\].RFW.BIT\[30\].FF REGF\[23\].RFW.CG\[3\]/GCLK DW[30] VGND VGND VPWR VPWR
+ REGF\[23\].RFW.BIT\[30\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[31\].RFW.BIT\[15\].OBUF2 REGF\[31\].RFW.BIT\[15\].FF/Q REGF\[31\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[15] sky130_fd_sc_hd__ebufn_2
Xfill_49_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_32_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[4\].RFW.BIT\[31\].OBUF1 REGF\[4\].RFW.BIT\[31\].FF/Q REGF\[4\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[31] sky130_fd_sc_hd__ebufn_2
Xfill_25_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.BIT\[18\].OBUF1 REGF\[3\].RFW.BIT\[18\].FF/Q REGF\[3\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[18] sky130_fd_sc_hd__ebufn_2
Xfill_18_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[16\].RFW.BIT\[24\].OBUF1 REGF\[16\].RFW.BIT\[24\].FF/Q REGF\[16\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[24] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.BIT\[11\].OBUF2 REGF\[29\].RFW.BIT\[11\].FF/Q REGF\[29\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[11] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.BIT\[13\].OBUF1 REGF\[21\].RFW.BIT\[13\].FF/Q REGF\[21\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[13] sky130_fd_sc_hd__ebufn_2
XREGF\[1\].RFW.BIT\[19\].FF REGF\[1\].RFW.CG\[2\]/GCLK DW[19] VGND VGND VPWR VPWR
+ REGF\[1\].RFW.BIT\[19\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[2\].RFW.CG\[3\] CLK REGF\[2\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[2\].RFW.CG\[3\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[7\].RFW.BIT\[13\].FF REGF\[7\].RFW.CG\[1\]/GCLK DW[13] VGND VGND VPWR VPWR
+ REGF\[7\].RFW.BIT\[13\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_29_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[22\].RFW.BIT\[29\].OBUF2 REGF\[22\].RFW.BIT\[29\].FF/Q REGF\[22\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[29] sky130_fd_sc_hd__ebufn_2
Xfill_45_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_45_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[7\].RFW.BIT\[19\].OBUF2 REGF\[7\].RFW.BIT\[19\].FF/Q REGF\[7\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[19] sky130_fd_sc_hd__ebufn_2
Xfill_61_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_22_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_61_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_61_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[28\].RFW.CG\[2\] CLK REGF\[28\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[28\].RFW.CG\[2\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_59_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.BIT\[27\].OBUF1 REGF\[12\].RFW.BIT\[27\].FF/Q REGF\[12\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[27] sky130_fd_sc_hd__ebufn_2
XREGF\[25\].RFW.BIT\[14\].OBUF2 REGF\[25\].RFW.BIT\[14\].FF/Q REGF\[25\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[14] sky130_fd_sc_hd__ebufn_2
Xfill_10_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_10_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_10_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[1\].RFW.CG\[0\] CLK REGF\[1\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[1\].RFW.CG\[0\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XDEC1.D2.ABUF\[1\] RB[1] VGND VGND VPWR VPWR DEC1.D2.AND7/B sky130_fd_sc_hd__clkbuf_2
XREGF\[24\].RFW.BIT\[13\].FF REGF\[24\].RFW.CG\[1\]/GCLK DW[13] VGND VGND VPWR VPWR
+ REGF\[24\].RFW.BIT\[13\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_19_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_19_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_19_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[15\].RFW.BIT\[12\].OBUF1 REGF\[15\].RFW.BIT\[12\].FF/Q REGF\[15\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[12] sky130_fd_sc_hd__ebufn_2
Xfill_35_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[31\].RFW.BIT\[3\].OBUF2 REGF\[31\].RFW.BIT\[3\].FF/Q REGF\[31\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[3] sky130_fd_sc_hd__ebufn_2
Xfill_51_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_51_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[30\].RFW.CGAND DEC2.D3.AND6/X WE VGND VGND VPWR VPWR REGF\[30\].RFW.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xgenblk1.RFW0.BIT\[28\].OBUF1 genblk1.RFW0.TIE\[3\]/LO genblk1.RFW0.INV1\[3\]/Y VGND
+ VGND VPWR VPWR DA[28] sky130_fd_sc_hd__ebufn_2
XREGF\[13\].RFW.BIT\[26\].FF REGF\[13\].RFW.CG\[3\]/GCLK DW[26] VGND VGND VPWR VPWR
+ REGF\[13\].RFW.BIT\[26\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_7_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XREGF\[16\].RFW.INV1\[0\] DEC0.D2.AND0/Y VGND VGND VPWR VPWR REGF\[16\].RFW.INV1\[0\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_7_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_7_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_7_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_7_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[16\].RFW.BIT\[28\].OBUF2 REGF\[16\].RFW.BIT\[28\].FF/Q REGF\[16\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[28] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.BIT\[20\].FF REGF\[19\].RFW.CG\[2\]/GCLK DW[20] VGND VGND VPWR VPWR
+ REGF\[19\].RFW.BIT\[20\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[21\].RFW.BIT\[17\].OBUF2 REGF\[21\].RFW.BIT\[17\].FF/Q REGF\[21\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[17] sky130_fd_sc_hd__ebufn_2
XREGF\[22\].RFW.BIT\[30\].OBUF2 REGF\[22\].RFW.BIT\[30\].FF/Q REGF\[22\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[30] sky130_fd_sc_hd__ebufn_2
Xfill_30_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_23_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[7\].RFW.BIT\[20\].OBUF2 REGF\[7\].RFW.BIT\[20\].FF/Q REGF\[7\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[20] sky130_fd_sc_hd__ebufn_2
Xfill_16_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.INV2\[1\] DEC1.D3.AND7/X VGND VGND VPWR VPWR REGF\[31\].RFW.INV2\[1\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[19\].RFW.BIT\[13\].OBUF2 REGF\[19\].RFW.BIT\[13\].FF/Q REGF\[19\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[13] sky130_fd_sc_hd__ebufn_2
Xtap_52_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[11\].RFW.BIT\[15\].OBUF1 REGF\[11\].RFW.BIT\[15\].FF/Q REGF\[11\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[15] sky130_fd_sc_hd__ebufn_2
Xtap_38_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_56_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_56_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_56_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[16\].RFW.CG\[2\] CLK REGF\[16\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[16\].RFW.CG\[2\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XDEC2.D3.AND2 DEC2.D3.AND7/C DEC2.D3.AND7/A DEC2.D3.AND7/B DEC2.D3.AND7/D VGND VGND
+ VPWR VPWR DEC2.D3.AND2/X sky130_fd_sc_hd__and4bb_2
Xfill_21_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_21_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.BIT\[23\].OBUF2 REGF\[3\].RFW.BIT\[23\].FF/Q REGF\[3\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[23] sky130_fd_sc_hd__ebufn_2
Xfill_21_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XREGF\[15\].RFW.BIT\[16\].OBUF2 REGF\[15\].RFW.BIT\[16\].FF/Q REGF\[15\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[16] sky130_fd_sc_hd__ebufn_2
XREGF\[8\].RFW.BIT\[19\].FF REGF\[8\].RFW.CG\[2\]/GCLK DW[19] VGND VGND VPWR VPWR
+ REGF\[8\].RFW.BIT\[19\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[10\].RFW.BIT\[11\].FF REGF\[10\].RFW.CG\[1\]/GCLK DW[11] VGND VGND VPWR VPWR
+ REGF\[10\].RFW.BIT\[11\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[4\].RFW.BIT\[21\].FF REGF\[4\].RFW.CG\[2\]/GCLK DW[21] VGND VGND VPWR VPWR
+ REGF\[4\].RFW.BIT\[21\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_7_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[10\].RFW.INV2\[1\] DEC1.D1.AND2/X VGND VGND VPWR VPWR REGF\[10\].RFW.INV2\[1\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[19\].RFW.BIT\[4\].FF REGF\[19\].RFW.CG\[0\]/GCLK DW[4] VGND VGND VPWR VPWR
+ REGF\[19\].RFW.BIT\[4\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[25\].RFW.BIT\[19\].FF REGF\[25\].RFW.CG\[2\]/GCLK DW[19] VGND VGND VPWR VPWR
+ REGF\[25\].RFW.BIT\[19\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_0_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[21\].RFW.BIT\[21\].FF REGF\[21\].RFW.CG\[2\]/GCLK DW[21] VGND VGND VPWR VPWR
+ REGF\[21\].RFW.BIT\[21\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[26\].RFW.INV2\[2\] DEC1.D3.AND2/X VGND VGND VPWR VPWR REGF\[26\].RFW.INV2\[2\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[11\].RFW.BIT\[19\].OBUF2 REGF\[11\].RFW.BIT\[19\].FF/Q REGF\[11\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[19] sky130_fd_sc_hd__ebufn_2
Xfill_42_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.BIT\[6\].FF REGF\[18\].RFW.CG\[0\]/GCLK DW[6] VGND VGND VPWR VPWR
+ REGF\[18\].RFW.BIT\[6\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[2\].RFW.BIT\[11\].OBUF2 REGF\[2\].RFW.BIT\[11\].FF/Q REGF\[2\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[11] sky130_fd_sc_hd__ebufn_2
Xtap_50_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_36_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[27\].RFW.BIT\[29\].OBUF1 REGF\[27\].RFW.BIT\[29\].FF/Q REGF\[27\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[29] sky130_fd_sc_hd__ebufn_2
Xtap_28_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_16_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[17\].RFW.BIT\[8\].FF REGF\[17\].RFW.CG\[1\]/GCLK DW[8] VGND VGND VPWR VPWR
+ REGF\[17\].RFW.BIT\[8\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_16_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC0.D3.ABUF\[2\] RA[2] VGND VGND VPWR VPWR DEC0.D3.AND7/C sky130_fd_sc_hd__clkbuf_2
Xfill_32_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_32_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[22\].RFW.INV1\[3\] DEC0.D2.AND6/X VGND VGND VPWR VPWR REGF\[22\].RFW.INV1\[3\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_57_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgenblk1.RFW0.INV1\[1\] DEC0.D0.AND0/Y VGND VGND VPWR VPWR genblk1.RFW0.INV1\[1\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_4_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_4_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_57_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[11\].RFW.BIT\[20\].OBUF2 REGF\[11\].RFW.BIT\[20\].FF/Q REGF\[11\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[20] sky130_fd_sc_hd__ebufn_2
Xfill_4_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_5_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[30\].RFW.BIT\[1\].OBUF2 REGF\[30\].RFW.BIT\[1\].FF/Q REGF\[30\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[1] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[17\].OBUF1 REGF\[26\].RFW.BIT\[17\].FF/Q REGF\[26\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[17] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[30\].OBUF1 REGF\[27\].RFW.BIT\[30\].FF/Q REGF\[27\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[30] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[27\].FF REGF\[5\].RFW.CG\[3\]/GCLK DW[27] VGND VGND VPWR VPWR
+ REGF\[5\].RFW.BIT\[27\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[11\].RFW.BIT\[17\].FF REGF\[11\].RFW.CG\[2\]/GCLK DW[17] VGND VGND VPWR VPWR
+ REGF\[11\].RFW.BIT\[17\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[17\].RFW.BIT\[11\].FF REGF\[17\].RFW.CG\[1\]/GCLK DW[11] VGND VGND VPWR VPWR
+ REGF\[17\].RFW.BIT\[11\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_37_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_53_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_53_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDEC2.D0.AND5 DEC2.D0.AND7/B DEC2.D0.AND7/A DEC2.D0.AND7/C DEC2.D0.AND7/D VGND VGND
+ VPWR VPWR DEC2.D0.AND5/X sky130_fd_sc_hd__and4b_2
Xtap_30_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_41_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[22\].RFW.BIT\[27\].FF REGF\[22\].RFW.CG\[3\]/GCLK DW[27] VGND VGND VPWR VPWR
+ REGF\[22\].RFW.BIT\[27\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_27_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[28\].RFW.BIT\[21\].FF REGF\[28\].RFW.CG\[2\]/GCLK DW[21] VGND VGND VPWR VPWR
+ REGF\[28\].RFW.BIT\[21\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_27_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_27_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[8\].RFW.BIT\[23\].OBUF1 REGF\[8\].RFW.BIT\[23\].FF/Q REGF\[8\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[23] sky130_fd_sc_hd__ebufn_2
Xfill_43_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_43_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_43_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_62_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_55_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC1.D1.AND7 DEC1.D1.AND7/A DEC1.D1.AND7/B DEC1.D1.AND7/C DEC1.D1.AND7/D VGND VGND
+ VPWR VPWR DEC1.D1.AND7/X sky130_fd_sc_hd__and4_2
Xfill_48_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[2\].RFW.BIT\[12\].FF REGF\[2\].RFW.CG\[1\]/GCLK DW[12] VGND VGND VPWR VPWR
+ REGF\[2\].RFW.BIT\[12\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_3_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[4\].RFW.BIT\[26\].OBUF1 REGF\[4\].RFW.BIT\[26\].FF/Q REGF\[4\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[26] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[19\].OBUF1 REGF\[16\].RFW.BIT\[19\].FF/Q REGF\[16\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[19] sky130_fd_sc_hd__ebufn_2
Xtap_20_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_48_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[22\].RFW.BIT\[21\].OBUF1 REGF\[22\].RFW.BIT\[21\].FF/Q REGF\[22\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[21] sky130_fd_sc_hd__ebufn_2
Xtap_6_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[7\].RFW.BIT\[11\].OBUF1 REGF\[7\].RFW.BIT\[11\].FF/Q REGF\[7\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[11] sky130_fd_sc_hd__ebufn_2
Xfill_13_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_13_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_13_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_13_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_13_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[8\].RFW.BIT\[27\].OBUF2 REGF\[8\].RFW.BIT\[27\].FF/Q REGF\[8\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[27] sky130_fd_sc_hd__ebufn_2
XREGF\[8\].RFW.INV2\[1\] DEC1.D1.AND0/Y VGND VGND VPWR VPWR REGF\[8\].RFW.INV2\[1\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[18\].RFW.BIT\[17\].FF REGF\[18\].RFW.CG\[2\]/GCLK DW[17] VGND VGND VPWR VPWR
+ REGF\[18\].RFW.BIT\[17\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_38_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_34_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_27_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[26\].RFW.BIT\[22\].OBUF2 REGF\[26\].RFW.BIT\[22\].FF/Q REGF\[26\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[22] sky130_fd_sc_hd__ebufn_2
XREGF\[30\].RFW.BIT\[22\].FF REGF\[30\].RFW.CG\[2\]/GCLK DW[22] VGND VGND VPWR VPWR
+ REGF\[30\].RFW.BIT\[22\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_1_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_1_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_1_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.BIT\[11\].OBUF2 REGF\[31\].RFW.BIT\[11\].FF/Q REGF\[31\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[11] sky130_fd_sc_hd__ebufn_2
XREGF\[3\].RFW.BIT\[14\].OBUF1 REGF\[3\].RFW.BIT\[14\].FF/Q REGF\[3\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[14] sky130_fd_sc_hd__ebufn_2
Xfill_60_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[16\].RFW.BIT\[20\].OBUF1 REGF\[16\].RFW.BIT\[20\].FF/Q REGF\[16\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[20] sky130_fd_sc_hd__ebufn_2
Xfill_53_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[29\].RFW.BIT\[27\].FF REGF\[29\].RFW.CG\[3\]/GCLK DW[27] VGND VGND VPWR VPWR
+ REGF\[29\].RFW.BIT\[27\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_46_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[24\].RFW.CG\[1\] CLK REGF\[24\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[24\].RFW.CG\[1\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[22\].RFW.BIT\[25\].OBUF2 REGF\[22\].RFW.BIT\[25\].FF/Q REGF\[22\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[25] sky130_fd_sc_hd__ebufn_2
Xfill_50_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[4\].RFW.INV1\[2\] DEC0.D0.AND4/X VGND VGND VPWR VPWR REGF\[4\].RFW.INV1\[2\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_59_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_59_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_59_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[7\].RFW.BIT\[15\].OBUF2 REGF\[7\].RFW.BIT\[15\].FF/Q REGF\[7\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[15] sky130_fd_sc_hd__ebufn_2
Xtap_11_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_36_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.BIT\[18\].FF REGF\[3\].RFW.CG\[2\]/GCLK DW[18] VGND VGND VPWR VPWR
+ REGF\[3\].RFW.BIT\[18\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_4_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.BIT\[23\].OBUF1 REGF\[12\].RFW.BIT\[23\].FF/Q REGF\[12\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[23] sky130_fd_sc_hd__ebufn_2
XREGF\[25\].RFW.BIT\[10\].OBUF2 REGF\[25\].RFW.BIT\[10\].FF/Q REGF\[25\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[10] sky130_fd_sc_hd__ebufn_2
XREGF\[9\].RFW.BIT\[12\].FF REGF\[9\].RFW.CG\[1\]/GCLK DW[12] VGND VGND VPWR VPWR
+ REGF\[9\].RFW.BIT\[12\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_24_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_24_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[24\].RFW.INV1\[0\] DEC0.D3.AND0/Y VGND VGND VPWR VPWR REGF\[24\].RFW.INV1\[0\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_40_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_40_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[14\].RFW.BIT\[1\].FF REGF\[14\].RFW.CG\[0\]/GCLK DW[1] VGND VGND VPWR VPWR
+ REGF\[14\].RFW.BIT\[1\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_49_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_49_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[18\].FF REGF\[20\].RFW.CG\[2\]/GCLK DW[18] VGND VGND VPWR VPWR
+ REGF\[20\].RFW.BIT\[18\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_32_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[4\].RFW.BIT\[31\].OBUF2 REGF\[4\].RFW.BIT\[31\].FF/Q REGF\[4\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[31] sky130_fd_sc_hd__ebufn_2
Xgenblk1.RFW0.BIT\[24\].OBUF1 genblk1.RFW0.TIE\[3\]/LO genblk1.RFW0.INV1\[3\]/Y VGND
+ VGND VPWR VPWR DA[24] sky130_fd_sc_hd__ebufn_2
Xfill_25_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.BIT\[18\].OBUF2 REGF\[3\].RFW.BIT\[18\].FF/Q REGF\[3\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[18] sky130_fd_sc_hd__ebufn_2
Xfill_18_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[16\].RFW.BIT\[24\].OBUF2 REGF\[16\].RFW.BIT\[24\].FF/Q REGF\[16\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[24] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[12\].FF REGF\[26\].RFW.CG\[1\]/GCLK DW[12] VGND VGND VPWR VPWR
+ REGF\[26\].RFW.BIT\[12\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[13\].RFW.BIT\[3\].FF REGF\[13\].RFW.CG\[0\]/GCLK DW[3] VGND VGND VPWR VPWR
+ REGF\[13\].RFW.BIT\[3\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[21\].RFW.BIT\[13\].OBUF2 REGF\[21\].RFW.BIT\[13\].FF/Q REGF\[21\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[13] sky130_fd_sc_hd__ebufn_2
XREGF\[12\].RFW.CG\[1\] CLK REGF\[12\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[12\].RFW.CG\[1\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[11\].RFW.BIT\[11\].OBUF1 REGF\[11\].RFW.BIT\[11\].FF/Q REGF\[11\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[11] sky130_fd_sc_hd__ebufn_2
XREGF\[15\].RFW.BIT\[25\].FF REGF\[15\].RFW.CG\[3\]/GCLK DW[25] VGND VGND VPWR VPWR
+ REGF\[15\].RFW.BIT\[25\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[12\].RFW.BIT\[5\].FF REGF\[12\].RFW.CG\[0\]/GCLK DW[5] VGND VGND VPWR VPWR
+ REGF\[12\].RFW.BIT\[5\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_45_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.BIT\[28\].FF REGF\[31\].RFW.CG\[3\]/GCLK DW[28] VGND VGND VPWR VPWR
+ REGF\[31\].RFW.BIT\[28\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_22_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_61_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_61_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_59_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.BIT\[27\].OBUF2 REGF\[12\].RFW.BIT\[27\].FF/Q REGF\[12\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[27] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[1\].FF REGF\[27\].RFW.CG\[0\]/GCLK DW[1] VGND VGND VPWR VPWR
+ REGF\[27\].RFW.BIT\[1\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_10_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_10_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_10_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[11\].RFW.BIT\[7\].FF REGF\[11\].RFW.CG\[0\]/GCLK DW[7] VGND VGND VPWR VPWR
+ REGF\[11\].RFW.BIT\[7\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_19_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_19_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_19_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XDEC2.D3.ENBUF DEC2.D.AND3/X VGND VGND VPWR VPWR DEC2.D3.AND7/D sky130_fd_sc_hd__clkbuf_2
XREGF\[19\].RFW.INV1\[1\] DEC0.D2.AND3/X VGND VGND VPWR VPWR REGF\[19\].RFW.INV1\[1\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[15\].RFW.BIT\[12\].OBUF2 REGF\[15\].RFW.BIT\[12\].FF/Q REGF\[15\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[12] sky130_fd_sc_hd__ebufn_2
Xfill_35_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_35_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[26\].RFW.BIT\[3\].FF REGF\[26\].RFW.CG\[0\]/GCLK DW[3] VGND VGND VPWR VPWR
+ REGF\[26\].RFW.BIT\[3\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[10\].RFW.BIT\[9\].FF REGF\[10\].RFW.CG\[1\]/GCLK DW[9] VGND VGND VPWR VPWR
+ REGF\[10\].RFW.BIT\[9\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_51_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_51_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_51_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgenblk1.RFW0.BIT\[28\].OBUF2 genblk1.RFW0.TIE\[7\]/LO genblk1.RFW0.INV2\[3\]/Y VGND
+ VGND VPWR VPWR DB[28] sky130_fd_sc_hd__ebufn_2
Xfill_7_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_7_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_7_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_7_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[25\].RFW.BIT\[5\].FF REGF\[25\].RFW.CG\[0\]/GCLK DW[5] VGND VGND VPWR VPWR
+ REGF\[25\].RFW.BIT\[5\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_30_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_23_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XREGF\[6\].RFW.BIT\[20\].FF REGF\[6\].RFW.CG\[2\]/GCLK DW[20] VGND VGND VPWR VPWR
+ REGF\[6\].RFW.BIT\[20\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[12\].RFW.BIT\[10\].FF REGF\[12\].RFW.CG\[1\]/GCLK DW[10] VGND VGND VPWR VPWR
+ REGF\[12\].RFW.BIT\[10\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_16_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDEC1.D0.ABUF\[0\] RB[0] VGND VGND VPWR VPWR DEC1.D0.AND7/A sky130_fd_sc_hd__clkbuf_2
XREGF\[11\].RFW.BIT\[15\].OBUF2 REGF\[11\].RFW.BIT\[15\].FF/Q REGF\[11\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[15] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[7\].FF REGF\[24\].RFW.CG\[0\]/GCLK DW[7] VGND VGND VPWR VPWR
+ REGF\[24\].RFW.BIT\[7\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_38_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_56_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[27\].RFW.BIT\[18\].FF REGF\[27\].RFW.CG\[2\]/GCLK DW[18] VGND VGND VPWR VPWR
+ REGF\[27\].RFW.BIT\[18\].FF/Q sky130_fd_sc_hd__dfxtp_1
XDEC2.D3.AND3 DEC2.D3.AND7/C DEC2.D3.AND7/B DEC2.D3.AND7/A DEC2.D3.AND7/D VGND VGND
+ VPWR VPWR DEC2.D3.AND3/X sky130_fd_sc_hd__and4b_2
XREGF\[23\].RFW.BIT\[20\].FF REGF\[23\].RFW.CG\[2\]/GCLK DW[20] VGND VGND VPWR VPWR
+ REGF\[23\].RFW.BIT\[20\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[27\].RFW.BIT\[25\].OBUF1 REGF\[27\].RFW.BIT\[25\].FF/Q REGF\[27\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[25] sky130_fd_sc_hd__ebufn_2
XREGF\[23\].RFW.BIT\[9\].FF REGF\[23\].RFW.CG\[1\]/GCLK DW[9] VGND VGND VPWR VPWR
+ REGF\[23\].RFW.BIT\[9\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[30\].RFW.INV1\[3\] DEC0.D3.AND6/X VGND VGND VPWR VPWR REGF\[30\].RFW.INV1\[3\]/Y
+ sky130_fd_sc_hd__inv_4
Xtap_57_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_21_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_21_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_21_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[9\].RFW.BIT\[4\].FF REGF\[9\].RFW.CG\[0\]/GCLK DW[4] VGND VGND VPWR VPWR REGF\[9\].RFW.BIT\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xfill_46_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[13\].RFW.INV2\[2\] DEC1.D1.AND5/X VGND VGND VPWR VPWR REGF\[13\].RFW.INV2\[2\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[29\].RFW.INV2\[3\] DEC1.D3.AND5/X VGND VGND VPWR VPWR REGF\[29\].RFW.INV2\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[8\].RFW.BIT\[6\].FF REGF\[8\].RFW.CG\[0\]/GCLK DW[6] VGND VGND VPWR VPWR REGF\[8\].RFW.BIT\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[23\].RFW.BIT\[28\].OBUF1 REGF\[23\].RFW.BIT\[28\].FF/Q REGF\[23\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[28] sky130_fd_sc_hd__ebufn_2
XREGF\[8\].RFW.BIT\[18\].OBUF1 REGF\[8\].RFW.BIT\[18\].FF/Q REGF\[8\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[18] sky130_fd_sc_hd__ebufn_2
XREGF\[9\].RFW.BIT\[31\].OBUF1 REGF\[9\].RFW.BIT\[31\].FF/Q REGF\[9\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[31] sky130_fd_sc_hd__ebufn_2
Xtap_0_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[26\].RFW.BIT\[13\].OBUF1 REGF\[26\].RFW.BIT\[13\].FF/Q REGF\[26\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[13] sky130_fd_sc_hd__ebufn_2
XREGF\[7\].RFW.BIT\[8\].FF REGF\[7\].RFW.CG\[1\]/GCLK DW[8] VGND VGND VPWR VPWR REGF\[7\].RFW.BIT\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xtap_50_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_36_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[27\].RFW.BIT\[29\].OBUF2 REGF\[27\].RFW.BIT\[29\].FF/Q REGF\[27\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[29] sky130_fd_sc_hd__ebufn_2
Xtap_28_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_44_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[7\].RFW.BIT\[26\].FF REGF\[7\].RFW.CG\[3\]/GCLK DW[26] VGND VGND VPWR VPWR
+ REGF\[7\].RFW.BIT\[26\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[13\].RFW.BIT\[16\].FF REGF\[13\].RFW.CG\[2\]/GCLK DW[16] VGND VGND VPWR VPWR
+ REGF\[13\].RFW.BIT\[16\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_16_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_16_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_16_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[17\].RFW.BIT\[27\].OBUF1 REGF\[17\].RFW.BIT\[27\].FF/Q REGF\[17\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[27] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.BIT\[10\].FF REGF\[19\].RFW.CG\[1\]/GCLK DW[10] VGND VGND VPWR VPWR
+ REGF\[19\].RFW.BIT\[10\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_32_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_32_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[22\].RFW.BIT\[16\].OBUF1 REGF\[22\].RFW.BIT\[16\].FF/Q REGF\[22\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[16] sky130_fd_sc_hd__ebufn_2
Xfill_57_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_4_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_4_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_57_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_57_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_4_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_5_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[24\].RFW.BIT\[26\].FF REGF\[24\].RFW.CG\[3\]/GCLK DW[26] VGND VGND VPWR VPWR
+ REGF\[24\].RFW.BIT\[26\].FF/Q sky130_fd_sc_hd__dfxtp_1
XDEC0.D1.ABUF\[1\] RA[1] VGND VGND VPWR VPWR DEC0.D1.AND7/B sky130_fd_sc_hd__clkbuf_2
XREGF\[26\].RFW.BIT\[17\].OBUF2 REGF\[26\].RFW.BIT\[17\].FF/Q REGF\[26\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[17] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[30\].OBUF2 REGF\[27\].RFW.BIT\[30\].FF/Q REGF\[27\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[30] sky130_fd_sc_hd__ebufn_2
Xtap_8_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[4\].RFW.BIT\[22\].OBUF1 REGF\[4\].RFW.BIT\[22\].FF/Q REGF\[4\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[22] sky130_fd_sc_hd__ebufn_2
Xfill_53_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[16\].RFW.BIT\[15\].OBUF1 REGF\[16\].RFW.BIT\[15\].FF/Q REGF\[16\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[15] sky130_fd_sc_hd__ebufn_2
XDEC2.D0.AND6 DEC2.D0.AND7/A DEC2.D0.AND7/B DEC2.D0.AND7/C DEC2.D0.AND7/D VGND VGND
+ VPWR VPWR DEC2.D0.AND6/X sky130_fd_sc_hd__and4b_2
Xtap_30_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[4\].RFW.BIT\[11\].FF REGF\[4\].RFW.CG\[1\]/GCLK DW[11] VGND VGND VPWR VPWR
+ REGF\[4\].RFW.BIT\[11\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_41_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_34_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[21\].RFW.CG\[3\] CLK REGF\[21\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[21\].RFW.CG\[3\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_27_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_27_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_27_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_27_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XREGF\[8\].RFW.BIT\[23\].OBUF2 REGF\[8\].RFW.BIT\[23\].FF/Q REGF\[8\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[23] sky130_fd_sc_hd__ebufn_2
Xfill_43_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_43_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_43_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_43_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[21\].RFW.BIT\[11\].FF REGF\[21\].RFW.CG\[1\]/GCLK DW[11] VGND VGND VPWR VPWR
+ REGF\[21\].RFW.BIT\[11\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[12\].RFW.BIT\[18\].OBUF1 REGF\[12\].RFW.BIT\[18\].FF/Q REGF\[12\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[18] sky130_fd_sc_hd__ebufn_2
XREGF\[13\].RFW.BIT\[31\].OBUF1 REGF\[13\].RFW.BIT\[31\].FF/Q REGF\[13\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[31] sky130_fd_sc_hd__ebufn_2
Xfill_62_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfill_55_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_48_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[9\].RFW.CG\[0\] CLK REGF\[9\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[9\].RFW.CG\[0\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[20\].RFW.CG\[0\] CLK REGF\[20\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[20\].RFW.CG\[0\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[3\].RFW.BIT\[10\].OBUF1 REGF\[3\].RFW.BIT\[10\].FF/Q REGF\[3\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[10] sky130_fd_sc_hd__ebufn_2
Xfill_3_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[10\].RFW.BIT\[24\].FF REGF\[10\].RFW.CG\[3\]/GCLK DW[24] VGND VGND VPWR VPWR
+ REGF\[10\].RFW.BIT\[24\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xgenblk1.RFW0.BIT\[19\].OBUF1 genblk1.RFW0.TIE\[2\]/LO genblk1.RFW0.INV1\[2\]/Y VGND
+ VGND VPWR VPWR DA[19] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.BIT\[26\].OBUF2 REGF\[4\].RFW.BIT\[26\].FF/Q REGF\[4\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[26] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[19\].OBUF2 REGF\[16\].RFW.BIT\[19\].FF/Q REGF\[16\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[19] sky130_fd_sc_hd__ebufn_2
Xtap_20_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_48_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[22\].RFW.BIT\[21\].OBUF2 REGF\[22\].RFW.BIT\[21\].FF/Q REGF\[22\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[21] sky130_fd_sc_hd__ebufn_2
Xtap_6_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[21\].RFW.BIT\[0\].FF REGF\[21\].RFW.CG\[0\]/GCLK DW[0] VGND VGND VPWR VPWR
+ REGF\[21\].RFW.BIT\[0\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[7\].RFW.BIT\[11\].OBUF2 REGF\[7\].RFW.BIT\[11\].FF/Q REGF\[7\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[11] sky130_fd_sc_hd__ebufn_2
Xfill_13_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_13_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_13_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_13_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[20\].RFW.BIT\[2\].FF REGF\[20\].RFW.CG\[0\]/GCLK DW[2] VGND VGND VPWR VPWR
+ REGF\[20\].RFW.BIT\[2\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_38_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_38_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_27_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_54_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_1_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_1_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[5\].RFW.BIT\[17\].FF REGF\[5\].RFW.CG\[2\]/GCLK DW[17] VGND VGND VPWR VPWR
+ REGF\[5\].RFW.BIT\[17\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xgenblk1.RFW0.BIT\[20\].OBUF1 genblk1.RFW0.TIE\[2\]/LO genblk1.RFW0.INV1\[2\]/Y VGND
+ VGND VPWR VPWR DA[20] sky130_fd_sc_hd__ebufn_2
XREGF\[3\].RFW.BIT\[14\].OBUF2 REGF\[3\].RFW.BIT\[14\].FF/Q REGF\[3\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[14] sky130_fd_sc_hd__ebufn_2
Xfill_60_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[16\].RFW.BIT\[20\].OBUF2 REGF\[16\].RFW.BIT\[20\].FF/Q REGF\[16\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[20] sky130_fd_sc_hd__ebufn_2
Xfill_53_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[7\].RFW.INV1\[3\] DEC0.D0.AND7/X VGND VGND VPWR VPWR REGF\[7\].RFW.INV1\[3\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_46_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_39_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[22\].RFW.BIT\[17\].FF REGF\[22\].RFW.CG\[2\]/GCLK DW[17] VGND VGND VPWR VPWR
+ REGF\[22\].RFW.BIT\[17\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[11\].RFW.INV1\[0\] DEC0.D1.AND3/X VGND VGND VPWR VPWR REGF\[11\].RFW.INV1\[0\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[28\].RFW.BIT\[11\].FF REGF\[28\].RFW.CG\[1\]/GCLK DW[11] VGND VGND VPWR VPWR
+ REGF\[28\].RFW.BIT\[11\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_59_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_59_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[27\].RFW.INV1\[1\] DEC0.D3.AND3/X VGND VGND VPWR VPWR REGF\[27\].RFW.INV1\[1\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[4\].RFW.BIT\[1\].FF REGF\[4\].RFW.CG\[0\]/GCLK DW[1] VGND VGND VPWR VPWR REGF\[4\].RFW.BIT\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xtap_11_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_36_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.BIT\[23\].OBUF2 REGF\[12\].RFW.BIT\[23\].FF/Q REGF\[12\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[23] sky130_fd_sc_hd__ebufn_2
Xtap_52_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_24_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_24_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_24_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[17\].RFW.BIT\[24\].FF REGF\[17\].RFW.CG\[3\]/GCLK DW[24] VGND VGND VPWR VPWR
+ REGF\[17\].RFW.BIT\[24\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[3\].RFW.BIT\[3\].FF REGF\[3\].RFW.CG\[0\]/GCLK DW[3] VGND VGND VPWR VPWR REGF\[3\].RFW.BIT\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xfill_40_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_40_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_49_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_49_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_49_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_32_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgenblk1.RFW0.BIT\[24\].OBUF2 genblk1.RFW0.TIE\[7\]/LO genblk1.RFW0.INV2\[3\]/Y VGND
+ VGND VPWR VPWR DB[24] sky130_fd_sc_hd__ebufn_2
Xfill_25_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.BIT\[6\].FF REGF\[31\].RFW.CG\[0\]/GCLK DW[6] VGND VGND VPWR VPWR
+ REGF\[31\].RFW.BIT\[6\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[2\].RFW.BIT\[5\].FF REGF\[2\].RFW.CG\[0\]/GCLK DW[5] VGND VGND VPWR VPWR REGF\[2\].RFW.BIT\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xfill_18_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[30\].RFW.BIT\[8\].FF REGF\[30\].RFW.CG\[1\]/GCLK DW[8] VGND VGND VPWR VPWR
+ REGF\[30\].RFW.BIT\[8\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[1\].RFW.BIT\[7\].FF REGF\[1\].RFW.CG\[0\]/GCLK DW[7] VGND VGND VPWR VPWR REGF\[1\].RFW.BIT\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[11\].RFW.BIT\[11\].OBUF2 REGF\[11\].RFW.BIT\[11\].FF/Q REGF\[11\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[11] sky130_fd_sc_hd__ebufn_2
Xfill_61_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[2\].RFW.BIT\[25\].FF REGF\[2\].RFW.CG\[3\]/GCLK DW[25] VGND VGND VPWR VPWR
+ REGF\[2\].RFW.BIT\[25\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[9\].RFW.BIT\[26\].OBUF1 REGF\[9\].RFW.BIT\[26\].FF/Q REGF\[9\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[26] sky130_fd_sc_hd__ebufn_2
Xfill_10_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[30\].RFW.BIT\[12\].FF REGF\[30\].RFW.CG\[1\]/GCLK DW[12] VGND VGND VPWR VPWR
+ REGF\[30\].RFW.BIT\[12\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_10_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_10_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[27\].RFW.BIT\[21\].OBUF1 REGF\[27\].RFW.BIT\[21\].FF/Q REGF\[27\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[21] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.INV2\[2\] DEC1.D2.AND5/X VGND VGND VPWR VPWR REGF\[21\].RFW.INV2\[2\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_19_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_19_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_19_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_19_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_19_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_51_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_51_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_51_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_51_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[29\].RFW.BIT\[17\].FF REGF\[29\].RFW.CG\[2\]/GCLK DW[17] VGND VGND VPWR VPWR
+ REGF\[29\].RFW.BIT\[17\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_7_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_7_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_7_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[5\].RFW.BIT\[29\].OBUF1 REGF\[5\].RFW.BIT\[29\].FF/Q REGF\[5\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[29] sky130_fd_sc_hd__ebufn_2
Xfill_7_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_7_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_30_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[23\].RFW.BIT\[24\].OBUF1 REGF\[23\].RFW.BIT\[24\].FF/Q REGF\[23\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[24] sky130_fd_sc_hd__ebufn_2
Xfill_23_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_16_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[8\].RFW.BIT\[14\].OBUF1 REGF\[8\].RFW.BIT\[14\].FF/Q REGF\[8\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[14] sky130_fd_sc_hd__ebufn_2
Xtap_38_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_56_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[27\].RFW.BIT\[25\].OBUF2 REGF\[27\].RFW.BIT\[25\].FF/Q REGF\[27\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[25] sky130_fd_sc_hd__ebufn_2
XDEC2.D3.AND4 DEC2.D3.AND7/A DEC2.D3.AND7/B DEC2.D3.AND7/C DEC2.D3.AND7/D VGND VGND
+ VPWR VPWR DEC2.D3.AND4/X sky130_fd_sc_hd__and4bb_2
Xtap_57_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[16\].RFW.INV2\[3\] DEC1.D2.AND0/Y VGND VGND VPWR VPWR REGF\[16\].RFW.INV2\[3\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_21_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[4\].RFW.BIT\[17\].OBUF1 REGF\[4\].RFW.BIT\[17\].FF/Q REGF\[4\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[17] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[30\].OBUF1 REGF\[5\].RFW.BIT\[30\].FF/Q REGF\[5\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[30] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.BIT\[23\].OBUF1 REGF\[17\].RFW.BIT\[23\].FF/Q REGF\[17\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[23] sky130_fd_sc_hd__ebufn_2
XREGF\[22\].RFW.BIT\[12\].OBUF1 REGF\[22\].RFW.BIT\[12\].FF/Q REGF\[22\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[12] sky130_fd_sc_hd__ebufn_2
Xfill_46_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_46_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_62_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[9\].RFW.BIT\[25\].FF REGF\[9\].RFW.CG\[3\]/GCLK DW[25] VGND VGND VPWR VPWR
+ REGF\[9\].RFW.BIT\[25\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[15\].RFW.BIT\[15\].FF REGF\[15\].RFW.CG\[1\]/GCLK DW[15] VGND VGND VPWR VPWR
+ REGF\[15\].RFW.BIT\[15\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[23\].RFW.BIT\[28\].OBUF2 REGF\[23\].RFW.BIT\[28\].FF/Q REGF\[23\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[28] sky130_fd_sc_hd__ebufn_2
XREGF\[31\].RFW.BIT\[18\].FF REGF\[31\].RFW.CG\[2\]/GCLK DW[18] VGND VGND VPWR VPWR
+ REGF\[31\].RFW.BIT\[18\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[9\].RFW.INV1\[0\] DEC0.D1.AND1/X VGND VGND VPWR VPWR REGF\[9\].RFW.INV1\[0\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[9\].RFW.BIT\[31\].OBUF2 REGF\[9\].RFW.BIT\[31\].FF/Q REGF\[9\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[31] sky130_fd_sc_hd__ebufn_2
XREGF\[8\].RFW.BIT\[18\].OBUF2 REGF\[8\].RFW.BIT\[18\].FF/Q REGF\[8\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[18] sky130_fd_sc_hd__ebufn_2
Xtap_0_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[13\].RFW.BIT\[26\].OBUF1 REGF\[13\].RFW.BIT\[26\].FF/Q REGF\[13\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[26] sky130_fd_sc_hd__ebufn_2
Xfill_21_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[26\].RFW.BIT\[13\].OBUF2 REGF\[26\].RFW.BIT\[13\].FF/Q REGF\[26\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[13] sky130_fd_sc_hd__ebufn_2
XDEC2.D2.ENBUF DEC2.D.AND2/X VGND VGND VPWR VPWR DEC2.D2.AND7/D sky130_fd_sc_hd__clkbuf_2
XREGF\[26\].RFW.BIT\[25\].FF REGF\[26\].RFW.CG\[3\]/GCLK DW[25] VGND VGND VPWR VPWR
+ REGF\[26\].RFW.BIT\[25\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_50_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_36_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.CG\[2\] CLK REGF\[6\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[6\].RFW.CG\[2\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[16\].RFW.BIT\[11\].OBUF1 REGF\[16\].RFW.BIT\[11\].FF/Q REGF\[16\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[11] sky130_fd_sc_hd__ebufn_2
Xtap_28_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_29_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_44_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_16_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_16_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_16_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_60_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[17\].RFW.BIT\[27\].OBUF2 REGF\[17\].RFW.BIT\[27\].FF/Q REGF\[17\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[27] sky130_fd_sc_hd__ebufn_2
Xfill_32_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_32_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_32_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[22\].RFW.BIT\[16\].OBUF2 REGF\[22\].RFW.BIT\[16\].FF/Q REGF\[22\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[16] sky130_fd_sc_hd__ebufn_2
XREGF\[6\].RFW.BIT\[10\].FF REGF\[6\].RFW.CG\[1\]/GCLK DW[10] VGND VGND VPWR VPWR
+ REGF\[6\].RFW.BIT\[10\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_57_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_4_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_57_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_57_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_57_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_4_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_4_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[12\].RFW.BIT\[14\].OBUF1 REGF\[12\].RFW.BIT\[14\].FF/Q REGF\[12\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[14] sky130_fd_sc_hd__ebufn_2
Xfill_5_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[3\].RFW.INV2\[1\] DEC1.D0.AND3/X VGND VGND VPWR VPWR REGF\[3\].RFW.INV2\[1\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[23\].RFW.BIT\[10\].FF REGF\[23\].RFW.CG\[1\]/GCLK DW[10] VGND VGND VPWR VPWR
+ REGF\[23\].RFW.BIT\[10\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xgenblk1.RFW0.BIT\[15\].OBUF1 genblk1.RFW0.TIE\[1\]/LO genblk1.RFW0.INV1\[1\]/Y VGND
+ VGND VPWR VPWR DA[15] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.BIT\[22\].OBUF2 REGF\[4\].RFW.BIT\[22\].FF/Q REGF\[4\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[22] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[15\].OBUF2 REGF\[16\].RFW.BIT\[15\].FF/Q REGF\[16\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[15] sky130_fd_sc_hd__ebufn_2
XDEC2.D0.AND7 DEC2.D0.AND7/A DEC2.D0.AND7/B DEC2.D0.AND7/C DEC2.D0.AND7/D VGND VGND
+ VPWR VPWR DEC2.D0.AND7/X sky130_fd_sc_hd__and4_2
XREGF\[12\].RFW.BIT\[23\].FF REGF\[12\].RFW.CG\[2\]/GCLK DW[23] VGND VGND VPWR VPWR
+ REGF\[12\].RFW.BIT\[23\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_34_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[2\].RFW.BIT\[9\].OBUF1 REGF\[2\].RFW.BIT\[9\].FF/Q REGF\[2\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[9] sky130_fd_sc_hd__ebufn_2
Xfill_27_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_27_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_27_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_27_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_27_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_43_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_43_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_43_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_43_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_43_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.BIT\[18\].OBUF2 REGF\[12\].RFW.BIT\[18\].FF/Q REGF\[12\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[18] sky130_fd_sc_hd__ebufn_2
XREGF\[13\].RFW.BIT\[31\].OBUF2 REGF\[13\].RFW.BIT\[31\].FF/Q REGF\[13\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[31] sky130_fd_sc_hd__ebufn_2
Xfill_62_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_55_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_48_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[3\].RFW.BIT\[10\].OBUF2 REGF\[3\].RFW.BIT\[10\].FF/Q REGF\[3\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[10] sky130_fd_sc_hd__ebufn_2
Xfill_3_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[28\].RFW.BIT\[28\].OBUF1 REGF\[28\].RFW.BIT\[28\].FF/Q REGF\[28\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[28] sky130_fd_sc_hd__ebufn_2
Xgenblk1.RFW0.BIT\[19\].OBUF2 genblk1.RFW0.TIE\[6\]/LO genblk1.RFW0.INV2\[2\]/Y VGND
+ VGND VPWR VPWR DB[19] sky130_fd_sc_hd__ebufn_2
XREGF\[7\].RFW.BIT\[16\].FF REGF\[7\].RFW.CG\[2\]/GCLK DW[16] VGND VGND VPWR VPWR
+ REGF\[7\].RFW.BIT\[16\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[4\].RFW.BIT\[9\].OBUF1 REGF\[4\].RFW.BIT\[9\].FF/Q REGF\[4\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[9] sky130_fd_sc_hd__ebufn_2
Xtap_20_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_6_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.INV2\[0\] DEC1.D2.AND2/X VGND VGND VPWR VPWR REGF\[18\].RFW.INV2\[0\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_13_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_13_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_13_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_13_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_13_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[24\].RFW.BIT\[16\].FF REGF\[24\].RFW.CG\[2\]/GCLK DW[16] VGND VGND VPWR VPWR
+ REGF\[24\].RFW.BIT\[16\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_38_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_38_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_54_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_54_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_1_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_1_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_1_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[27\].RFW.BIT\[16\].OBUF1 REGF\[27\].RFW.BIT\[16\].FF/Q REGF\[27\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[16] sky130_fd_sc_hd__ebufn_2
XREGF\[6\].RFW.BIT\[9\].OBUF1 REGF\[6\].RFW.BIT\[9\].FF/Q REGF\[6\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[9] sky130_fd_sc_hd__ebufn_2
XREGF\[13\].RFW.BIT\[29\].FF REGF\[13\].RFW.CG\[3\]/GCLK DW[29] VGND VGND VPWR VPWR
+ REGF\[13\].RFW.BIT\[29\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xgenblk1.RFW0.BIT\[20\].OBUF2 genblk1.RFW0.TIE\[6\]/LO genblk1.RFW0.INV2\[2\]/Y VGND
+ VGND VPWR VPWR DB[20] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.BIT\[23\].FF REGF\[19\].RFW.CG\[2\]/GCLK DW[23] VGND VGND VPWR VPWR
+ REGF\[19\].RFW.BIT\[23\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_60_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_53_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_46_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[14\].RFW.INV1\[1\] DEC0.D1.AND6/X VGND VGND VPWR VPWR REGF\[14\].RFW.INV1\[1\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_39_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_1_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDEC0.D1.AND0 DEC0.D1.AND7/A DEC0.D1.AND7/B DEC0.D1.AND7/C DEC0.D1.AND7/D VGND VGND
+ VPWR VPWR DEC0.D1.AND0/Y sky130_fd_sc_hd__nor4b_2
XREGF\[23\].RFW.BIT\[19\].OBUF1 REGF\[23\].RFW.BIT\[19\].FF/Q REGF\[23\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[19] sky130_fd_sc_hd__ebufn_2
Xfill_59_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[9\].RFW.BIT\[22\].OBUF1 REGF\[9\].RFW.BIT\[22\].FF/Q REGF\[9\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[22] sky130_fd_sc_hd__ebufn_2
Xtap_11_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_36_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[8\].RFW.BIT\[9\].OBUF1 REGF\[8\].RFW.BIT\[9\].FF/Q REGF\[8\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[9] sky130_fd_sc_hd__ebufn_2
Xtap_4_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_52_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_24_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_24_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_24_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[11\].RFW.BIT\[8\].OBUF1 REGF\[11\].RFW.BIT\[8\].FF/Q REGF\[11\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[8] sky130_fd_sc_hd__ebufn_2
Xfill_40_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_40_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_40_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[10\].RFW.BIT\[14\].FF REGF\[10\].RFW.CG\[1\]/GCLK DW[14] VGND VGND VPWR VPWR
+ REGF\[10\].RFW.BIT\[14\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[4\].RFW.BIT\[24\].FF REGF\[4\].RFW.CG\[3\]/GCLK DW[24] VGND VGND VPWR VPWR
+ REGF\[4\].RFW.BIT\[24\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_49_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_49_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_49_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_49_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[1\].RFW.BIT\[7\].OBUF1 REGF\[1\].RFW.BIT\[7\].FF/Q REGF\[1\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[7] sky130_fd_sc_hd__ebufn_2
Xfill_32_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_25_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[5\].RFW.BIT\[25\].OBUF1 REGF\[5\].RFW.BIT\[25\].FF/Q REGF\[5\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[25] sky130_fd_sc_hd__ebufn_2
Xfill_18_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[17\].RFW.BIT\[18\].OBUF1 REGF\[17\].RFW.BIT\[18\].FF/Q REGF\[17\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[18] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.BIT\[31\].OBUF1 REGF\[18\].RFW.BIT\[31\].FF/Q REGF\[18\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[31] sky130_fd_sc_hd__ebufn_2
XREGF\[23\].RFW.BIT\[20\].OBUF1 REGF\[23\].RFW.BIT\[20\].FF/Q REGF\[23\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[20] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.BIT\[7\].FF REGF\[19\].RFW.CG\[0\]/GCLK DW[7] VGND VGND VPWR VPWR
+ REGF\[19\].RFW.BIT\[7\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[21\].RFW.BIT\[24\].FF REGF\[21\].RFW.CG\[3\]/GCLK DW[24] VGND VGND VPWR VPWR
+ REGF\[21\].RFW.BIT\[24\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[8\].RFW.BIT\[10\].OBUF1 REGF\[8\].RFW.BIT\[10\].FF/Q REGF\[8\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[10] sky130_fd_sc_hd__ebufn_2
Xfill_51_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[13\].RFW.BIT\[8\].OBUF1 REGF\[13\].RFW.BIT\[8\].FF/Q REGF\[13\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[8] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.INV2\[3\] DEC1.D3.AND0/Y VGND VGND VPWR VPWR REGF\[24\].RFW.INV2\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[18\].RFW.BIT\[9\].FF REGF\[18\].RFW.CG\[1\]/GCLK DW[9] VGND VGND VPWR VPWR
+ REGF\[18\].RFW.BIT\[9\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[9\].RFW.BIT\[26\].OBUF2 REGF\[9\].RFW.BIT\[26\].FF/Q REGF\[9\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[26] sky130_fd_sc_hd__ebufn_2
XREGF\[1\].RFW.BIT\[28\].OBUF1 REGF\[1\].RFW.BIT\[28\].FF/Q REGF\[1\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[28] sky130_fd_sc_hd__ebufn_2
Xfill_10_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[3\].RFW.BIT\[7\].OBUF1 REGF\[3\].RFW.BIT\[7\].FF/Q REGF\[3\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[7] sky130_fd_sc_hd__ebufn_2
Xfill_10_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_10_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[27\].RFW.BIT\[21\].OBUF2 REGF\[27\].RFW.BIT\[21\].FF/Q REGF\[27\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[21] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[31\].FF REGF\[16\].RFW.CG\[3\]/GCLK DW[31] VGND VGND VPWR VPWR
+ REGF\[16\].RFW.BIT\[31\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_19_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_19_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_19_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_19_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xtap_2_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[4\].RFW.BIT\[13\].OBUF1 REGF\[4\].RFW.BIT\[13\].FF/Q REGF\[4\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[13] sky130_fd_sc_hd__ebufn_2
Xfill_35_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_35_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_35_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_51_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_51_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_51_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_51_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_51_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_7_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_7_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_7_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[5\].RFW.BIT\[29\].OBUF2 REGF\[5\].RFW.BIT\[29\].FF/Q REGF\[5\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[29] sky130_fd_sc_hd__ebufn_2
Xfill_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_7_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[15\].RFW.BIT\[8\].OBUF1 REGF\[15\].RFW.BIT\[8\].FF/Q REGF\[15\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[8] sky130_fd_sc_hd__ebufn_2
Xfill_30_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[23\].RFW.BIT\[24\].OBUF2 REGF\[23\].RFW.BIT\[24\].FF/Q REGF\[23\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[24] sky130_fd_sc_hd__ebufn_2
Xfill_23_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_16_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[29\].RFW.CG\[3\] CLK REGF\[29\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[29\].RFW.CG\[3\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[8\].RFW.BIT\[14\].OBUF2 REGF\[8\].RFW.BIT\[14\].FF/Q REGF\[8\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[14] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[7\].OBUF1 REGF\[5\].RFW.BIT\[7\].FF/Q REGF\[5\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[7] sky130_fd_sc_hd__ebufn_2
XREGF\[2\].RFW.CG\[1\] CLK REGF\[2\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[2\].RFW.CG\[1\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[13\].RFW.BIT\[22\].OBUF1 REGF\[13\].RFW.BIT\[22\].FF/Q REGF\[13\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[22] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.BIT\[14\].FF REGF\[17\].RFW.CG\[1\]/GCLK DW[14] VGND VGND VPWR VPWR
+ REGF\[17\].RFW.BIT\[14\].FF/Q sky130_fd_sc_hd__dfxtp_1
XDEC2.D3.AND5 DEC2.D3.AND7/B DEC2.D3.AND7/A DEC2.D3.AND7/C DEC2.D3.AND7/D VGND VGND
+ VPWR VPWR DEC2.D3.AND5/X sky130_fd_sc_hd__and4b_2
XREGF\[28\].RFW.CG\[0\] CLK REGF\[28\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[28\].RFW.CG\[0\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[17\].RFW.BIT\[8\].OBUF1 REGF\[17\].RFW.BIT\[8\].FF/Q REGF\[17\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[8] sky130_fd_sc_hd__ebufn_2
Xtap_57_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_21_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_21_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_21_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_58_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[4\].RFW.BIT\[17\].OBUF2 REGF\[4\].RFW.BIT\[17\].FF/Q REGF\[4\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[17] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[30\].OBUF2 REGF\[5\].RFW.BIT\[30\].FF/Q REGF\[5\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[30] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.BIT\[23\].OBUF2 REGF\[17\].RFW.BIT\[23\].FF/Q REGF\[17\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[23] sky130_fd_sc_hd__ebufn_2
XREGF\[7\].RFW.BIT\[7\].OBUF1 REGF\[7\].RFW.BIT\[7\].FF/Q REGF\[7\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[7] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.BIT\[24\].FF REGF\[28\].RFW.CG\[3\]/GCLK DW[24] VGND VGND VPWR VPWR
+ REGF\[28\].RFW.BIT\[24\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[22\].RFW.BIT\[12\].OBUF2 REGF\[22\].RFW.BIT\[12\].FF/Q REGF\[22\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[12] sky130_fd_sc_hd__ebufn_2
Xfill_46_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_46_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_62_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[10\].RFW.BIT\[6\].OBUF1 REGF\[10\].RFW.BIT\[6\].FF/Q REGF\[10\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[6] sky130_fd_sc_hd__ebufn_2
XREGF\[12\].RFW.BIT\[10\].OBUF1 REGF\[12\].RFW.BIT\[10\].FF/Q REGF\[12\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[10] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.CG\[3\] CLK REGF\[17\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[17\].RFW.CG\[3\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[2\].RFW.BIT\[15\].FF REGF\[2\].RFW.CG\[1\]/GCLK DW[15] VGND VGND VPWR VPWR
+ REGF\[2\].RFW.BIT\[15\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[19\].RFW.BIT\[8\].OBUF1 REGF\[19\].RFW.BIT\[8\].FF/Q REGF\[19\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[8] sky130_fd_sc_hd__ebufn_2
XREGF\[13\].RFW.BIT\[26\].OBUF2 REGF\[13\].RFW.BIT\[26\].FF/Q REGF\[13\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[26] sky130_fd_sc_hd__ebufn_2
Xfill_21_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_14_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgenblk1.RFW0.BIT\[11\].OBUF1 genblk1.RFW0.TIE\[1\]/LO genblk1.RFW0.INV1\[1\]/Y VGND
+ VGND VPWR VPWR DA[11] sky130_fd_sc_hd__ebufn_2
Xtap_50_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[9\].RFW.BIT\[7\].OBUF1 REGF\[9\].RFW.BIT\[7\].FF/Q REGF\[9\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[7] sky130_fd_sc_hd__ebufn_2
Xtap_36_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[16\].RFW.BIT\[11\].OBUF2 REGF\[16\].RFW.BIT\[11\].FF/Q REGF\[16\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[11] sky130_fd_sc_hd__ebufn_2
XREGF\[12\].RFW.BIT\[6\].OBUF1 REGF\[12\].RFW.BIT\[6\].FF/Q REGF\[12\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[6] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.CG\[0\] CLK REGF\[16\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[16\].RFW.CG\[0\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_44_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_16_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_16_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_16_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xtap_60_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_32_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_32_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_62_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_32_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[2\].RFW.BIT\[5\].OBUF1 REGF\[2\].RFW.BIT\[5\].FF/Q REGF\[2\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[5] sky130_fd_sc_hd__ebufn_2
Xfill_4_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_57_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_57_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_57_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_57_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[14\].RFW.BIT\[22\].FF REGF\[14\].RFW.CG\[2\]/GCLK DW[22] VGND VGND VPWR VPWR
+ REGF\[14\].RFW.BIT\[22\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_4_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_4_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[30\].RFW.BIT\[25\].FF REGF\[30\].RFW.CG\[3\]/GCLK DW[25] VGND VGND VPWR VPWR
+ REGF\[30\].RFW.BIT\[25\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[12\].RFW.BIT\[14\].OBUF2 REGF\[12\].RFW.BIT\[14\].FF/Q REGF\[12\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[14] sky130_fd_sc_hd__ebufn_2
XREGF\[6\].RFW.INV2\[2\] DEC1.D0.AND6/X VGND VGND VPWR VPWR REGF\[6\].RFW.INV2\[2\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_5_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[30\].RFW.BIT\[28\].OBUF1 REGF\[30\].RFW.BIT\[28\].FF/Q REGF\[30\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[28] sky130_fd_sc_hd__ebufn_2
XREGF\[14\].RFW.BIT\[6\].OBUF1 REGF\[14\].RFW.BIT\[6\].FF/Q REGF\[14\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[6] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.BIT\[24\].OBUF1 REGF\[28\].RFW.BIT\[24\].FF/Q REGF\[28\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[24] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.INV2\[0\] DEC1.D3.AND2/X VGND VGND VPWR VPWR REGF\[26\].RFW.INV2\[0\]/Y
+ sky130_fd_sc_hd__inv_4
Xgenblk1.RFW0.BIT\[15\].OBUF2 genblk1.RFW0.TIE\[5\]/LO genblk1.RFW0.INV2\[1\]/Y VGND
+ VGND VPWR VPWR DB[15] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[0\].FF REGF\[16\].RFW.CG\[0\]/GCLK DW[0] VGND VGND VPWR VPWR
+ REGF\[16\].RFW.BIT\[0\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[4\].RFW.BIT\[5\].OBUF1 REGF\[4\].RFW.BIT\[5\].FF/Q REGF\[4\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[5] sky130_fd_sc_hd__ebufn_2
Xtap_34_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[15\].RFW.BIT\[2\].FF REGF\[15\].RFW.CG\[0\]/GCLK DW[2] VGND VGND VPWR VPWR
+ REGF\[15\].RFW.BIT\[2\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[2\].RFW.INV1\[3\] DEC0.D0.AND2/X VGND VGND VPWR VPWR REGF\[2\].RFW.INV1\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[2\].RFW.BIT\[9\].OBUF2 REGF\[2\].RFW.BIT\[9\].FF/Q REGF\[2\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[9] sky130_fd_sc_hd__ebufn_2
Xfill_27_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[9\].RFW.BIT\[15\].FF REGF\[9\].RFW.CG\[1\]/GCLK DW[15] VGND VGND VPWR VPWR
+ REGF\[9\].RFW.BIT\[15\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_27_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_27_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_27_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[24\].RFW.BIT\[27\].OBUF1 REGF\[24\].RFW.BIT\[27\].FF/Q REGF\[24\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[27] sky130_fd_sc_hd__ebufn_2
XDEC0.D3.ABUF\[0\] RA[0] VGND VGND VPWR VPWR DEC0.D3.AND7/A sky130_fd_sc_hd__clkbuf_2
Xfill_43_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_43_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_43_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[16\].RFW.BIT\[6\].OBUF1 REGF\[16\].RFW.BIT\[6\].FF/Q REGF\[16\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[6] sky130_fd_sc_hd__ebufn_2
Xfill_43_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_43_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_43_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[9\].RFW.BIT\[17\].OBUF1 REGF\[9\].RFW.BIT\[17\].FF/Q REGF\[9\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[17] sky130_fd_sc_hd__ebufn_2
XREGF\[14\].RFW.BIT\[4\].FF REGF\[14\].RFW.CG\[0\]/GCLK DW[4] VGND VGND VPWR VPWR
+ REGF\[14\].RFW.BIT\[4\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[22\].RFW.INV1\[1\] DEC0.D2.AND6/X VGND VGND VPWR VPWR REGF\[22\].RFW.INV1\[1\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[27\].RFW.BIT\[12\].OBUF1 REGF\[27\].RFW.BIT\[12\].FF/Q REGF\[27\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[12] sky130_fd_sc_hd__ebufn_2
Xfill_62_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.BIT\[5\].OBUF1 REGF\[6\].RFW.BIT\[5\].FF/Q REGF\[6\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[5] sky130_fd_sc_hd__ebufn_2
Xfill_55_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_48_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XDEC2.D1.ENBUF DEC2.D.AND1/X VGND VGND VPWR VPWR DEC2.D1.AND7/D sky130_fd_sc_hd__clkbuf_2
XREGF\[29\].RFW.BIT\[0\].FF REGF\[29\].RFW.CG\[0\]/GCLK DW[0] VGND VGND VPWR VPWR
+ REGF\[29\].RFW.BIT\[0\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[26\].RFW.BIT\[15\].FF REGF\[26\].RFW.CG\[1\]/GCLK DW[15] VGND VGND VPWR VPWR
+ REGF\[26\].RFW.BIT\[15\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_3_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[13\].RFW.BIT\[6\].FF REGF\[13\].RFW.CG\[0\]/GCLK DW[6] VGND VGND VPWR VPWR
+ REGF\[13\].RFW.BIT\[6\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[28\].RFW.BIT\[28\].OBUF2 REGF\[28\].RFW.BIT\[28\].FF/Q REGF\[28\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[28] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.BIT\[9\].OBUF2 REGF\[4\].RFW.BIT\[9\].FF/Q REGF\[4\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[9] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.BIT\[2\].FF REGF\[28\].RFW.CG\[0\]/GCLK DW[2] VGND VGND VPWR VPWR
+ REGF\[28\].RFW.BIT\[2\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[12\].RFW.BIT\[8\].FF REGF\[12\].RFW.CG\[1\]/GCLK DW[8] VGND VGND VPWR VPWR
+ REGF\[12\].RFW.BIT\[8\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[15\].RFW.BIT\[28\].FF REGF\[15\].RFW.CG\[3\]/GCLK DW[28] VGND VGND VPWR VPWR
+ REGF\[15\].RFW.BIT\[28\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[18\].RFW.BIT\[26\].OBUF1 REGF\[18\].RFW.BIT\[26\].FF/Q REGF\[18\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[26] sky130_fd_sc_hd__ebufn_2
XREGF\[11\].RFW.BIT\[30\].FF REGF\[11\].RFW.CG\[3\]/GCLK DW[30] VGND VGND VPWR VPWR
+ REGF\[11\].RFW.BIT\[30\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[18\].RFW.BIT\[6\].OBUF1 REGF\[18\].RFW.BIT\[6\].FF/Q REGF\[18\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[6] sky130_fd_sc_hd__ebufn_2
Xtap_6_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[23\].RFW.BIT\[15\].OBUF1 REGF\[23\].RFW.BIT\[15\].FF/Q REGF\[23\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[15] sky130_fd_sc_hd__ebufn_2
Xfill_13_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_13_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_13_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_13_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[27\].RFW.BIT\[4\].FF REGF\[27\].RFW.CG\[0\]/GCLK DW[4] VGND VGND VPWR VPWR
+ REGF\[27\].RFW.BIT\[4\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[8\].RFW.BIT\[5\].OBUF1 REGF\[8\].RFW.BIT\[5\].FF/Q REGF\[8\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[5] sky130_fd_sc_hd__ebufn_2
Xtap_32_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[11\].RFW.BIT\[4\].OBUF1 REGF\[11\].RFW.BIT\[4\].FF/Q REGF\[11\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[4] sky130_fd_sc_hd__ebufn_2
Xfill_38_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_38_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_38_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[26\].RFW.BIT\[6\].FF REGF\[26\].RFW.CG\[0\]/GCLK DW[6] VGND VGND VPWR VPWR
+ REGF\[26\].RFW.BIT\[6\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_54_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_54_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[14\].RFW.BIT\[29\].OBUF1 REGF\[14\].RFW.BIT\[29\].FF/Q REGF\[14\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[29] sky130_fd_sc_hd__ebufn_2
Xfill_1_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[27\].RFW.BIT\[16\].OBUF2 REGF\[27\].RFW.BIT\[16\].FF/Q REGF\[27\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[16] sky130_fd_sc_hd__ebufn_2
XREGF\[6\].RFW.BIT\[9\].OBUF2 REGF\[6\].RFW.BIT\[9\].FF/Q REGF\[6\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[9] sky130_fd_sc_hd__ebufn_2
XREGF\[1\].RFW.BIT\[3\].OBUF1 REGF\[1\].RFW.BIT\[3\].FF/Q REGF\[1\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[3] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.INV1\[2\] DEC0.D2.AND1/X VGND VGND VPWR VPWR REGF\[17\].RFW.INV1\[2\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[20\].RFW.BIT\[31\].OBUF1 REGF\[20\].RFW.BIT\[31\].FF/Q REGF\[20\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[31] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[21\].OBUF1 REGF\[5\].RFW.BIT\[21\].FF/Q REGF\[5\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[21] sky130_fd_sc_hd__ebufn_2
Xfill_60_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[17\].RFW.BIT\[14\].OBUF1 REGF\[17\].RFW.BIT\[14\].FF/Q REGF\[17\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[14] sky130_fd_sc_hd__ebufn_2
XREGF\[25\].RFW.BIT\[8\].FF REGF\[25\].RFW.CG\[1\]/GCLK DW[8] VGND VGND VPWR VPWR
+ REGF\[25\].RFW.BIT\[8\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_53_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_46_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[6\].RFW.BIT\[23\].FF REGF\[6\].RFW.CG\[2\]/GCLK DW[23] VGND VGND VPWR VPWR
+ REGF\[6\].RFW.BIT\[23\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[12\].RFW.BIT\[13\].FF REGF\[12\].RFW.CG\[1\]/GCLK DW[13] VGND VGND VPWR VPWR
+ REGF\[12\].RFW.BIT\[13\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_1_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[13\].RFW.BIT\[4\].OBUF1 REGF\[13\].RFW.BIT\[4\].FF/Q REGF\[13\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[4] sky130_fd_sc_hd__ebufn_2
XDEC0.D1.AND1 DEC0.D1.AND7/C DEC0.D1.AND7/B DEC0.D1.AND7/A DEC0.D1.AND7/D VGND VGND
+ VPWR VPWR DEC0.D1.AND1/X sky130_fd_sc_hd__and4bb_2
XREGF\[23\].RFW.BIT\[19\].OBUF2 REGF\[23\].RFW.BIT\[19\].FF/Q REGF\[23\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[19] sky130_fd_sc_hd__ebufn_2
XREGF\[9\].RFW.BIT\[22\].OBUF2 REGF\[9\].RFW.BIT\[22\].FF/Q REGF\[9\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[22] sky130_fd_sc_hd__ebufn_2
XREGF\[8\].RFW.BIT\[9\].OBUF2 REGF\[8\].RFW.BIT\[9\].FF/Q REGF\[8\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[9] sky130_fd_sc_hd__ebufn_2
Xtap_4_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[1\].RFW.BIT\[24\].OBUF1 REGF\[1\].RFW.BIT\[24\].FF/Q REGF\[1\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[24] sky130_fd_sc_hd__ebufn_2
XREGF\[3\].RFW.BIT\[3\].OBUF1 REGF\[3\].RFW.BIT\[3\].FF/Q REGF\[3\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[3] sky130_fd_sc_hd__ebufn_2
Xtap_52_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[13\].RFW.BIT\[17\].OBUF1 REGF\[13\].RFW.BIT\[17\].FF/Q REGF\[13\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[17] sky130_fd_sc_hd__ebufn_2
XREGF\[23\].RFW.BIT\[23\].FF REGF\[23\].RFW.CG\[2\]/GCLK DW[23] VGND VGND VPWR VPWR
+ REGF\[23\].RFW.BIT\[23\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[14\].RFW.BIT\[30\].OBUF1 REGF\[14\].RFW.BIT\[30\].FF/Q REGF\[14\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[30] sky130_fd_sc_hd__ebufn_2
Xfill_24_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_24_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_24_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[11\].RFW.BIT\[8\].OBUF2 REGF\[11\].RFW.BIT\[8\].FF/Q REGF\[11\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[8] sky130_fd_sc_hd__ebufn_2
Xfill_40_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_40_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_40_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[9\].RFW.BIT\[7\].FF REGF\[9\].RFW.CG\[0\]/GCLK DW[7] VGND VGND VPWR VPWR REGF\[9\].RFW.BIT\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xfill_49_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_49_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_49_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_49_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_49_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[1\].RFW.BIT\[7\].OBUF2 REGF\[1\].RFW.BIT\[7\].FF/Q REGF\[1\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[7] sky130_fd_sc_hd__ebufn_2
Xfill_32_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[25\].RFW.CG\[2\] CLK REGF\[25\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[25\].RFW.CG\[2\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[18\].RFW.BIT\[30\].FF REGF\[18\].RFW.CG\[3\]/GCLK DW[30] VGND VGND VPWR VPWR
+ REGF\[18\].RFW.BIT\[30\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_25_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[5\].RFW.BIT\[25\].OBUF2 REGF\[5\].RFW.BIT\[25\].FF/Q REGF\[5\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[25] sky130_fd_sc_hd__ebufn_2
XREGF\[15\].RFW.BIT\[4\].OBUF1 REGF\[15\].RFW.BIT\[4\].FF/Q REGF\[15\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[4] sky130_fd_sc_hd__ebufn_2
Xfill_18_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[17\].RFW.BIT\[18\].OBUF2 REGF\[17\].RFW.BIT\[18\].FF/Q REGF\[17\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[18] sky130_fd_sc_hd__ebufn_2
XREGF\[8\].RFW.BIT\[9\].FF REGF\[8\].RFW.CG\[1\]/GCLK DW[9] VGND VGND VPWR VPWR REGF\[8\].RFW.BIT\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[18\].RFW.BIT\[31\].OBUF2 REGF\[18\].RFW.BIT\[31\].FF/Q REGF\[18\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[31] sky130_fd_sc_hd__ebufn_2
XREGF\[11\].RFW.INV2\[3\] DEC1.D1.AND3/X VGND VGND VPWR VPWR REGF\[11\].RFW.INV2\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[23\].RFW.BIT\[20\].OBUF2 REGF\[23\].RFW.BIT\[20\].FF/Q REGF\[23\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[20] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[3\].OBUF1 REGF\[5\].RFW.BIT\[3\].FF/Q REGF\[5\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[3] sky130_fd_sc_hd__ebufn_2
XREGF\[8\].RFW.BIT\[10\].OBUF2 REGF\[8\].RFW.BIT\[10\].FF/Q REGF\[8\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[10] sky130_fd_sc_hd__ebufn_2
Xfill_51_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_44_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[13\].RFW.BIT\[8\].OBUF2 REGF\[13\].RFW.BIT\[8\].FF/Q REGF\[13\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[8] sky130_fd_sc_hd__ebufn_2
XREGF\[1\].RFW.BIT\[28\].OBUF2 REGF\[1\].RFW.BIT\[28\].FF/Q REGF\[1\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[28] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.INV1\[0\] DEC0.D0.AND4/X VGND VGND VPWR VPWR REGF\[4\].RFW.INV1\[0\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[3\].RFW.BIT\[7\].OBUF2 REGF\[3\].RFW.BIT\[7\].FF/Q REGF\[3\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[7] sky130_fd_sc_hd__ebufn_2
Xfill_10_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_10_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_10_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[17\].RFW.BIT\[4\].OBUF1 REGF\[17\].RFW.BIT\[4\].FF/Q REGF\[17\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[4] sky130_fd_sc_hd__ebufn_2
Xfill_19_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_19_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_19_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_19_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_19_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[7\].RFW.BIT\[29\].FF REGF\[7\].RFW.CG\[3\]/GCLK DW[29] VGND VGND VPWR VPWR
+ REGF\[7\].RFW.BIT\[29\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[13\].RFW.BIT\[19\].FF REGF\[13\].RFW.CG\[2\]/GCLK DW[19] VGND VGND VPWR VPWR
+ REGF\[13\].RFW.BIT\[19\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xgenblk1.RFW0.BIT\[8\].OBUF1 genblk1.RFW0.TIE\[1\]/LO genblk1.RFW0.INV1\[1\]/Y VGND
+ VGND VPWR VPWR DA[8] sky130_fd_sc_hd__ebufn_2
Xtap_2_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.BIT\[31\].FF REGF\[3\].RFW.CG\[3\]/GCLK DW[31] VGND VGND VPWR VPWR
+ REGF\[3\].RFW.BIT\[31\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[4\].RFW.BIT\[13\].OBUF2 REGF\[4\].RFW.BIT\[13\].FF/Q REGF\[4\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[13] sky130_fd_sc_hd__ebufn_2
Xfill_35_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_35_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_35_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[19\].RFW.BIT\[13\].FF REGF\[19\].RFW.CG\[1\]/GCLK DW[13] VGND VGND VPWR VPWR
+ REGF\[19\].RFW.BIT\[13\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_35_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_51_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_51_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[7\].RFW.BIT\[3\].OBUF1 REGF\[7\].RFW.BIT\[3\].FF/Q REGF\[7\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[3] sky130_fd_sc_hd__ebufn_2
Xfill_51_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_51_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_51_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_51_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[13\].RFW.CG\[2\] CLK REGF\[13\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[13\].RFW.CG\[2\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_7_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_7_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_7_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_7_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_7_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[15\].RFW.BIT\[8\].OBUF2 REGF\[15\].RFW.BIT\[8\].FF/Q REGF\[15\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[8] sky130_fd_sc_hd__ebufn_2
XREGF\[10\].RFW.BIT\[2\].OBUF1 REGF\[10\].RFW.BIT\[2\].FF/Q REGF\[10\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[2] sky130_fd_sc_hd__ebufn_2
Xfill_30_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_23_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[24\].RFW.BIT\[29\].FF REGF\[24\].RFW.CG\[3\]/GCLK DW[29] VGND VGND VPWR VPWR
+ REGF\[24\].RFW.BIT\[29\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[20\].RFW.BIT\[31\].FF REGF\[20\].RFW.CG\[3\]/GCLK DW[31] VGND VGND VPWR VPWR
+ REGF\[20\].RFW.BIT\[31\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_16_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[5\].RFW.BIT\[7\].OBUF2 REGF\[5\].RFW.BIT\[7\].FF/Q REGF\[5\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[7] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.BIT\[4\].OBUF1 REGF\[19\].RFW.BIT\[4\].FF/Q REGF\[19\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[4] sky130_fd_sc_hd__ebufn_2
XREGF\[13\].RFW.BIT\[22\].OBUF2 REGF\[13\].RFW.BIT\[22\].FF/Q REGF\[13\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[22] sky130_fd_sc_hd__ebufn_2
XREGF\[9\].RFW.BIT\[3\].OBUF1 REGF\[9\].RFW.BIT\[3\].FF/Q REGF\[9\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[3] sky130_fd_sc_hd__ebufn_2
XDEC2.D3.AND6 DEC2.D3.AND7/A DEC2.D3.AND7/B DEC2.D3.AND7/C DEC2.D3.AND7/D VGND VGND
+ VPWR VPWR DEC2.D3.AND6/X sky130_fd_sc_hd__and4b_2
XREGF\[28\].RFW.BIT\[19\].OBUF1 REGF\[28\].RFW.BIT\[19\].FF/Q REGF\[28\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[19] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.BIT\[14\].FF REGF\[4\].RFW.CG\[1\]/GCLK DW[14] VGND VGND VPWR VPWR
+ REGF\[4\].RFW.BIT\[14\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[12\].RFW.BIT\[2\].OBUF1 REGF\[12\].RFW.BIT\[2\].FF/Q REGF\[12\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[2] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.BIT\[8\].OBUF2 REGF\[17\].RFW.BIT\[8\].FF/Q REGF\[17\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[8] sky130_fd_sc_hd__ebufn_2
Xtap_57_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_21_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_58_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[7\].RFW.BIT\[7\].OBUF2 REGF\[7\].RFW.BIT\[7\].FF/Q REGF\[7\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[7] sky130_fd_sc_hd__ebufn_2
XREGF\[2\].RFW.BIT\[1\].OBUF1 REGF\[2\].RFW.BIT\[1\].FF/Q REGF\[2\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[1] sky130_fd_sc_hd__ebufn_2
Xfill_46_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_46_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_46_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_62_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_62_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[10\].RFW.BIT\[6\].OBUF2 REGF\[10\].RFW.BIT\[6\].FF/Q REGF\[10\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[6] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.BIT\[14\].FF REGF\[21\].RFW.CG\[1\]/GCLK DW[14] VGND VGND VPWR VPWR
+ REGF\[21\].RFW.BIT\[14\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[12\].RFW.BIT\[10\].OBUF2 REGF\[12\].RFW.BIT\[10\].FF/Q REGF\[12\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[10] sky130_fd_sc_hd__ebufn_2
Xgenblk1.RFW0.TIE\[7\] VGND VGND VPWR VPWR genblk1.RFW0.TIE\[7\]/HI genblk1.RFW0.TIE\[7\]/LO
+ sky130_fd_sc_hd__conb_1
XREGF\[30\].RFW.BIT\[24\].OBUF1 REGF\[30\].RFW.BIT\[24\].FF/Q REGF\[30\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[24] sky130_fd_sc_hd__ebufn_2
XREGF\[14\].RFW.BIT\[2\].OBUF1 REGF\[14\].RFW.BIT\[2\].FF/Q REGF\[14\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[2] sky130_fd_sc_hd__ebufn_2
XREGF\[10\].RFW.BIT\[27\].FF REGF\[10\].RFW.CG\[3\]/GCLK DW[27] VGND VGND VPWR VPWR
+ REGF\[10\].RFW.BIT\[27\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_21_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XREGF\[19\].RFW.BIT\[8\].OBUF2 REGF\[19\].RFW.BIT\[8\].FF/Q REGF\[19\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[8] sky130_fd_sc_hd__ebufn_2
Xfill_14_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[28\].RFW.BIT\[20\].OBUF1 REGF\[28\].RFW.BIT\[20\].FF/Q REGF\[28\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[20] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[21\].FF REGF\[16\].RFW.CG\[2\]/GCLK DW[21] VGND VGND VPWR VPWR
+ REGF\[16\].RFW.BIT\[21\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[22\].RFW.BIT\[1\].FF REGF\[22\].RFW.CG\[0\]/GCLK DW[1] VGND VGND VPWR VPWR
+ REGF\[22\].RFW.BIT\[1\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[9\].RFW.BIT\[7\].OBUF2 REGF\[9\].RFW.BIT\[7\].FF/Q REGF\[9\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[7] sky130_fd_sc_hd__ebufn_2
Xgenblk1.RFW0.BIT\[11\].OBUF2 genblk1.RFW0.TIE\[5\]/LO genblk1.RFW0.INV2\[1\]/Y VGND
+ VGND VPWR VPWR DB[11] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.BIT\[1\].OBUF1 REGF\[4\].RFW.BIT\[1\].FF/Q REGF\[4\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[1] sky130_fd_sc_hd__ebufn_2
Xtap_36_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.BIT\[6\].OBUF2 REGF\[12\].RFW.BIT\[6\].FF/Q REGF\[12\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[6] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.BIT\[3\].FF REGF\[21\].RFW.CG\[0\]/GCLK DW[3] VGND VGND VPWR VPWR
+ REGF\[21\].RFW.BIT\[3\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_16_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_16_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_60_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.BIT\[28\].OBUF1 REGF\[6\].RFW.BIT\[28\].FF/Q REGF\[6\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[28] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[31\].FF REGF\[27\].RFW.CG\[3\]/GCLK DW[31] VGND VGND VPWR VPWR
+ REGF\[27\].RFW.BIT\[31\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_32_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_32_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_62_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_32_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[30\].RFW.INV1\[1\] DEC0.D3.AND6/X VGND VGND VPWR VPWR REGF\[30\].RFW.INV1\[1\]/Y
+ sky130_fd_sc_hd__inv_4
Xtap_55_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[2\].RFW.BIT\[5\].OBUF2 REGF\[2\].RFW.BIT\[5\].FF/Q REGF\[2\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[5] sky130_fd_sc_hd__ebufn_2
XREGF\[9\].RFW.INV2\[3\] DEC1.D1.AND1/X VGND VGND VPWR VPWR REGF\[9\].RFW.INV2\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[24\].RFW.BIT\[23\].OBUF1 REGF\[24\].RFW.BIT\[23\].FF/Q REGF\[24\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[23] sky130_fd_sc_hd__ebufn_2
XREGF\[20\].RFW.BIT\[5\].FF REGF\[20\].RFW.CG\[0\]/GCLK DW[5] VGND VGND VPWR VPWR
+ REGF\[20\].RFW.BIT\[5\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[16\].RFW.BIT\[2\].OBUF1 REGF\[16\].RFW.BIT\[2\].FF/Q REGF\[16\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[2] sky130_fd_sc_hd__ebufn_2
XREGF\[9\].RFW.BIT\[13\].OBUF1 REGF\[9\].RFW.BIT\[13\].FF/Q REGF\[9\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[13] sky130_fd_sc_hd__ebufn_2
Xfill_57_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_57_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_57_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_57_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_4_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfill_4_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_4_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_57_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[13\].RFW.INV2\[0\] DEC1.D1.AND5/X VGND VGND VPWR VPWR REGF\[13\].RFW.INV2\[0\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[6\].RFW.BIT\[0\].FF REGF\[6\].RFW.CG\[0\]/GCLK DW[0] VGND VGND VPWR VPWR REGF\[6\].RFW.BIT\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[1\].RFW.BIT\[22\].FF REGF\[1\].RFW.CG\[2\]/GCLK DW[22] VGND VGND VPWR VPWR
+ REGF\[1\].RFW.BIT\[22\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[6\].RFW.BIT\[1\].OBUF1 REGF\[6\].RFW.BIT\[1\].FF/Q REGF\[6\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[1] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.INV2\[1\] DEC1.D3.AND5/X VGND VGND VPWR VPWR REGF\[29\].RFW.INV2\[1\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[30\].RFW.BIT\[28\].OBUF2 REGF\[30\].RFW.BIT\[28\].FF/Q REGF\[30\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[28] sky130_fd_sc_hd__ebufn_2
XREGF\[14\].RFW.BIT\[6\].OBUF2 REGF\[14\].RFW.BIT\[6\].FF/Q REGF\[14\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[6] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.BIT\[24\].OBUF2 REGF\[28\].RFW.BIT\[24\].FF/Q REGF\[28\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[24] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[2\].FF REGF\[5\].RFW.CG\[0\]/GCLK DW[2] VGND VGND VPWR VPWR REGF\[5\].RFW.BIT\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[20\].RFW.BIT\[26\].OBUF1 REGF\[20\].RFW.BIT\[26\].FF/Q REGF\[20\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[26] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[16\].OBUF1 REGF\[5\].RFW.BIT\[16\].FF/Q REGF\[5\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[16] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.BIT\[5\].OBUF2 REGF\[4\].RFW.BIT\[5\].FF/Q REGF\[4\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[5] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.BIT\[22\].OBUF1 REGF\[18\].RFW.BIT\[22\].FF/Q REGF\[18\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[22] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.BIT\[2\].OBUF1 REGF\[18\].RFW.BIT\[2\].FF/Q REGF\[18\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[2] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.BIT\[14\].FF REGF\[28\].RFW.CG\[1\]/GCLK DW[14] VGND VGND VPWR VPWR
+ REGF\[28\].RFW.BIT\[14\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[23\].RFW.BIT\[11\].OBUF1 REGF\[23\].RFW.BIT\[11\].FF/Q REGF\[23\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[11] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.BIT\[4\].FF REGF\[4\].RFW.CG\[0\]/GCLK DW[4] VGND VGND VPWR VPWR REGF\[4\].RFW.BIT\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xtap_34_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_27_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_27_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[8\].RFW.BIT\[1\].OBUF1 REGF\[8\].RFW.BIT\[1\].FF/Q REGF\[8\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[1] sky130_fd_sc_hd__ebufn_2
Xfill_27_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_27_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_27_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_27_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[24\].RFW.BIT\[27\].OBUF2 REGF\[24\].RFW.BIT\[27\].FF/Q REGF\[24\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[27] sky130_fd_sc_hd__ebufn_2
XREGF\[25\].RFW.INV1\[2\] DEC0.D3.AND1/X VGND VGND VPWR VPWR REGF\[25\].RFW.INV1\[2\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[17\].RFW.BIT\[27\].FF REGF\[17\].RFW.CG\[3\]/GCLK DW[27] VGND VGND VPWR VPWR
+ REGF\[17\].RFW.BIT\[27\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_43_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_43_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_43_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[11\].RFW.BIT\[0\].OBUF1 REGF\[11\].RFW.BIT\[0\].FF/Q REGF\[11\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[0] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[6\].OBUF2 REGF\[16\].RFW.BIT\[6\].FF/Q REGF\[16\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[6] sky130_fd_sc_hd__ebufn_2
Xfill_43_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_43_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_43_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[3\].RFW.BIT\[6\].FF REGF\[3\].RFW.CG\[0\]/GCLK DW[6] VGND VGND VPWR VPWR REGF\[3\].RFW.BIT\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[9\].RFW.BIT\[17\].OBUF2 REGF\[9\].RFW.BIT\[17\].FF/Q REGF\[9\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[17] sky130_fd_sc_hd__ebufn_2
XREGF\[1\].RFW.BIT\[19\].OBUF1 REGF\[1\].RFW.BIT\[19\].FF/Q REGF\[1\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[19] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[12\].OBUF2 REGF\[27\].RFW.BIT\[12\].FF/Q REGF\[27\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[12] sky130_fd_sc_hd__ebufn_2
Xfill_62_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[14\].RFW.BIT\[25\].OBUF1 REGF\[14\].RFW.BIT\[25\].FF/Q REGF\[14\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[25] sky130_fd_sc_hd__ebufn_2
XREGF\[6\].RFW.BIT\[5\].OBUF2 REGF\[6\].RFW.BIT\[5\].FF/Q REGF\[6\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[5] sky130_fd_sc_hd__ebufn_2
Xfill_55_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_48_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[31\].RFW.BIT\[9\].FF REGF\[31\].RFW.CG\[1\]/GCLK DW[9] VGND VGND VPWR VPWR
+ REGF\[31\].RFW.BIT\[9\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[2\].RFW.BIT\[8\].FF REGF\[2\].RFW.CG\[1\]/GCLK DW[8] VGND VGND VPWR VPWR REGF\[2\].RFW.BIT\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xfill_3_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[17\].RFW.BIT\[10\].OBUF1 REGF\[17\].RFW.BIT\[10\].FF/Q REGF\[17\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[10] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.BIT\[26\].OBUF2 REGF\[18\].RFW.BIT\[26\].FF/Q REGF\[18\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[26] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.BIT\[6\].OBUF2 REGF\[18\].RFW.BIT\[6\].FF/Q REGF\[18\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[6] sky130_fd_sc_hd__ebufn_2
XREGF\[13\].RFW.BIT\[0\].OBUF1 REGF\[13\].RFW.BIT\[0\].FF/Q REGF\[13\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[0] sky130_fd_sc_hd__ebufn_2
Xtap_6_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[23\].RFW.BIT\[15\].OBUF2 REGF\[23\].RFW.BIT\[15\].FF/Q REGF\[23\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[15] sky130_fd_sc_hd__ebufn_2
XREGF\[10\].RFW.BIT\[28\].OBUF1 REGF\[10\].RFW.BIT\[28\].FF/Q REGF\[10\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[28] sky130_fd_sc_hd__ebufn_2
XREGF\[2\].RFW.BIT\[28\].FF REGF\[2\].RFW.CG\[3\]/GCLK DW[28] VGND VGND VPWR VPWR
+ REGF\[2\].RFW.BIT\[28\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_13_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_13_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[9\].OBUF1 REGF\[20\].RFW.BIT\[9\].FF/Q REGF\[20\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[9] sky130_fd_sc_hd__ebufn_2
XREGF\[8\].RFW.BIT\[22\].FF REGF\[8\].RFW.CG\[2\]/GCLK DW[22] VGND VGND VPWR VPWR
+ REGF\[8\].RFW.BIT\[22\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[14\].RFW.BIT\[12\].FF REGF\[14\].RFW.CG\[1\]/GCLK DW[12] VGND VGND VPWR VPWR
+ REGF\[14\].RFW.BIT\[12\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_13_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_13_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_13_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[8\].RFW.BIT\[5\].OBUF2 REGF\[8\].RFW.BIT\[5\].FF/Q REGF\[8\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[5] sky130_fd_sc_hd__ebufn_2
XREGF\[1\].RFW.BIT\[20\].OBUF1 REGF\[1\].RFW.BIT\[20\].FF/Q REGF\[1\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[20] sky130_fd_sc_hd__ebufn_2
XREGF\[30\].RFW.BIT\[15\].FF REGF\[30\].RFW.CG\[1\]/GCLK DW[15] VGND VGND VPWR VPWR
+ REGF\[30\].RFW.BIT\[15\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[13\].RFW.BIT\[13\].OBUF1 REGF\[13\].RFW.BIT\[13\].FF/Q REGF\[13\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[13] sky130_fd_sc_hd__ebufn_2
Xtap_32_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[11\].RFW.BIT\[4\].OBUF2 REGF\[11\].RFW.BIT\[4\].FF/Q REGF\[11\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[4] sky130_fd_sc_hd__ebufn_2
Xtap_18_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[21\].RFW.CG\[1\] CLK REGF\[21\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[21\].RFW.CG\[1\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_38_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_38_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_38_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC1.D0.AND0 DEC1.D0.AND7/A DEC1.D0.AND7/B DEC1.D0.AND7/C DEC1.D0.AND7/D VGND VGND
+ VPWR VPWR DEC1.D0.AND0/Y sky130_fd_sc_hd__nor4b_2
Xfill_54_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_54_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_54_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[14\].RFW.BIT\[29\].OBUF2 REGF\[14\].RFW.BIT\[29\].FF/Q REGF\[14\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[29] sky130_fd_sc_hd__ebufn_2
Xfill_1_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_1_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[1\].RFW.BIT\[3\].OBUF2 REGF\[1\].RFW.BIT\[3\].FF/Q REGF\[1\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[3] sky130_fd_sc_hd__ebufn_2
XREGF\[20\].RFW.BIT\[31\].OBUF2 REGF\[20\].RFW.BIT\[31\].FF/Q REGF\[20\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[31] sky130_fd_sc_hd__ebufn_2
XREGF\[25\].RFW.BIT\[22\].FF REGF\[25\].RFW.CG\[2\]/GCLK DW[22] VGND VGND VPWR VPWR
+ REGF\[25\].RFW.BIT\[22\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[5\].RFW.BIT\[21\].OBUF2 REGF\[5\].RFW.BIT\[21\].FF/Q REGF\[5\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[21] sky130_fd_sc_hd__ebufn_2
XREGF\[15\].RFW.BIT\[0\].OBUF1 REGF\[15\].RFW.BIT\[0\].FF/Q REGF\[15\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[0] sky130_fd_sc_hd__ebufn_2
Xfill_60_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_53_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[17\].RFW.BIT\[14\].OBUF2 REGF\[17\].RFW.BIT\[14\].FF/Q REGF\[17\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[14] sky130_fd_sc_hd__ebufn_2
Xfill_46_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[22\].RFW.BIT\[9\].OBUF1 REGF\[22\].RFW.BIT\[9\].FF/Q REGF\[22\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[9] sky130_fd_sc_hd__ebufn_2
Xfill_1_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC0.D1.AND2 DEC0.D1.AND7/C DEC0.D1.AND7/A DEC0.D1.AND7/B DEC0.D1.AND7/D VGND VGND
+ VPWR VPWR DEC0.D1.AND2/X sky130_fd_sc_hd__and4bb_2
XREGF\[13\].RFW.BIT\[4\].OBUF2 REGF\[13\].RFW.BIT\[4\].FF/Q REGF\[13\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[4] sky130_fd_sc_hd__ebufn_2
Xtap_4_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[1\].RFW.BIT\[24\].OBUF2 REGF\[1\].RFW.BIT\[24\].FF/Q REGF\[1\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[24] sky130_fd_sc_hd__ebufn_2
XREGF\[3\].RFW.BIT\[3\].OBUF2 REGF\[3\].RFW.BIT\[3\].FF/Q REGF\[3\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[3] sky130_fd_sc_hd__ebufn_2
XREGF\[14\].RFW.BIT\[30\].OBUF2 REGF\[14\].RFW.BIT\[30\].FF/Q REGF\[14\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[30] sky130_fd_sc_hd__ebufn_2
XREGF\[13\].RFW.BIT\[17\].OBUF2 REGF\[13\].RFW.BIT\[17\].FF/Q REGF\[13\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[17] sky130_fd_sc_hd__ebufn_2
Xfill_24_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_24_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_24_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[17\].RFW.BIT\[0\].OBUF1 REGF\[17\].RFW.BIT\[0\].FF/Q REGF\[17\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[0] sky130_fd_sc_hd__ebufn_2
Xfill_40_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgenblk1.RFW0.BIT\[4\].OBUF1 genblk1.RFW0.TIE\[0\]/LO genblk1.RFW0.INV1\[0\]/Y VGND
+ VGND VPWR VPWR DA[4] sky130_fd_sc_hd__ebufn_2
XDEC2.D0.ENBUF DEC2.D.AND0/Y VGND VGND VPWR VPWR DEC2.D0.AND7/D sky130_fd_sc_hd__clkbuf_2
Xfill_40_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_40_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[24\].RFW.BIT\[9\].OBUF1 REGF\[24\].RFW.BIT\[9\].FF/Q REGF\[24\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[9] sky130_fd_sc_hd__ebufn_2
Xfill_49_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_49_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[29\].RFW.BIT\[27\].OBUF1 REGF\[29\].RFW.BIT\[27\].FF/Q REGF\[29\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[27] sky130_fd_sc_hd__ebufn_2
Xfill_49_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_49_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_49_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_49_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_25_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_18_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[15\].RFW.BIT\[4\].OBUF2 REGF\[15\].RFW.BIT\[4\].FF/Q REGF\[15\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[4] sky130_fd_sc_hd__ebufn_2
XREGF\[9\].RFW.BIT\[28\].FF REGF\[9\].RFW.CG\[3\]/GCLK DW[28] VGND VGND VPWR VPWR
+ REGF\[9\].RFW.BIT\[28\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[15\].RFW.BIT\[18\].FF REGF\[15\].RFW.CG\[2\]/GCLK DW[18] VGND VGND VPWR VPWR
+ REGF\[15\].RFW.BIT\[18\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[5\].RFW.BIT\[30\].FF REGF\[5\].RFW.CG\[3\]/GCLK DW[30] VGND VGND VPWR VPWR
+ REGF\[5\].RFW.BIT\[30\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[11\].RFW.BIT\[20\].FF REGF\[11\].RFW.CG\[2\]/GCLK DW[20] VGND VGND VPWR VPWR
+ REGF\[11\].RFW.BIT\[20\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[5\].RFW.BIT\[3\].OBUF2 REGF\[5\].RFW.BIT\[3\].FF/Q REGF\[5\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[3] sky130_fd_sc_hd__ebufn_2
Xfill_51_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[7\].RFW.INV1\[1\] DEC0.D0.AND7/X VGND VGND VPWR VPWR REGF\[7\].RFW.INV1\[1\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_44_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_37_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[19\].RFW.BIT\[0\].OBUF1 REGF\[19\].RFW.BIT\[0\].FF/Q REGF\[19\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[0] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[9\].OBUF1 REGF\[26\].RFW.BIT\[9\].FF/Q REGF\[26\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[9] sky130_fd_sc_hd__ebufn_2
XREGF\[30\].RFW.BIT\[19\].OBUF1 REGF\[30\].RFW.BIT\[19\].FF/Q REGF\[30\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[19] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[28\].FF REGF\[26\].RFW.CG\[3\]/GCLK DW[28] VGND VGND VPWR VPWR
+ REGF\[26\].RFW.BIT\[28\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[22\].RFW.BIT\[30\].FF REGF\[22\].RFW.CG\[3\]/GCLK DW[30] VGND VGND VPWR VPWR
+ REGF\[22\].RFW.BIT\[30\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_10_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_10_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_10_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[28\].RFW.BIT\[15\].OBUF1 REGF\[28\].RFW.BIT\[15\].FF/Q REGF\[28\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[15] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.BIT\[4\].OBUF2 REGF\[17\].RFW.BIT\[4\].FF/Q REGF\[17\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[4] sky130_fd_sc_hd__ebufn_2
Xfill_19_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_19_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_19_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_19_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgenblk1.RFW0.BIT\[8\].OBUF2 genblk1.RFW0.TIE\[5\]/LO genblk1.RFW0.INV2\[1\]/Y VGND
+ VGND VPWR VPWR DB[8] sky130_fd_sc_hd__ebufn_2
Xtap_2_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_35_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_51_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_51_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[7\].RFW.BIT\[3\].OBUF2 REGF\[7\].RFW.BIT\[3\].FF/Q REGF\[7\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[3] sky130_fd_sc_hd__ebufn_2
Xfill_51_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_51_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_51_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_51_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[6\].RFW.BIT\[13\].FF REGF\[6\].RFW.CG\[1\]/GCLK DW[13] VGND VGND VPWR VPWR
+ REGF\[6\].RFW.BIT\[13\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_7_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_7_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_7_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_7_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_7_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[10\].RFW.BIT\[2\].OBUF2 REGF\[10\].RFW.BIT\[2\].FF/Q REGF\[10\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[2] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.BIT\[29\].OBUF1 REGF\[19\].RFW.BIT\[29\].FF/Q REGF\[19\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[29] sky130_fd_sc_hd__ebufn_2
Xfill_30_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[28\].RFW.BIT\[9\].OBUF1 REGF\[28\].RFW.BIT\[9\].FF/Q REGF\[28\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[9] sky130_fd_sc_hd__ebufn_2
Xfill_23_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[24\].RFW.BIT\[18\].OBUF1 REGF\[24\].RFW.BIT\[18\].FF/Q REGF\[24\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[18] sky130_fd_sc_hd__ebufn_2
XREGF\[25\].RFW.BIT\[31\].OBUF1 REGF\[25\].RFW.BIT\[31\].FF/Q REGF\[25\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[31] sky130_fd_sc_hd__ebufn_2
Xfill_16_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[30\].RFW.BIT\[20\].OBUF1 REGF\[30\].RFW.BIT\[20\].FF/Q REGF\[30\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[20] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.BIT\[4\].OBUF2 REGF\[19\].RFW.BIT\[4\].FF/Q REGF\[19\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[4] sky130_fd_sc_hd__ebufn_2
XREGF\[23\].RFW.BIT\[13\].FF REGF\[23\].RFW.CG\[1\]/GCLK DW[13] VGND VGND VPWR VPWR
+ REGF\[23\].RFW.BIT\[13\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[21\].RFW.BIT\[7\].OBUF1 REGF\[21\].RFW.BIT\[7\].FF/Q REGF\[21\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[7] sky130_fd_sc_hd__ebufn_2
XREGF\[1\].RFW.INV2\[2\] DEC1.D0.AND1/X VGND VGND VPWR VPWR REGF\[1\].RFW.INV2\[2\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[9\].RFW.BIT\[3\].OBUF2 REGF\[9\].RFW.BIT\[3\].FF/Q REGF\[9\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[3] sky130_fd_sc_hd__ebufn_2
XDEC2.D3.AND7 DEC2.D3.AND7/A DEC2.D3.AND7/B DEC2.D3.AND7/C DEC2.D3.AND7/D VGND VGND
+ VPWR VPWR DEC2.D3.AND7/X sky130_fd_sc_hd__and4_2
XREGF\[28\].RFW.BIT\[19\].OBUF2 REGF\[28\].RFW.BIT\[19\].FF/Q REGF\[28\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[19] sky130_fd_sc_hd__ebufn_2
XREGF\[12\].RFW.BIT\[26\].FF REGF\[12\].RFW.CG\[3\]/GCLK DW[26] VGND VGND VPWR VPWR
+ REGF\[12\].RFW.BIT\[26\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[12\].RFW.BIT\[2\].OBUF2 REGF\[12\].RFW.BIT\[2\].FF/Q REGF\[12\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[2] sky130_fd_sc_hd__ebufn_2
Xfill_21_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_21_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xtap_58_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.BIT\[20\].FF REGF\[18\].RFW.CG\[2\]/GCLK DW[20] VGND VGND VPWR VPWR
+ REGF\[18\].RFW.BIT\[20\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[6\].RFW.BIT\[24\].OBUF1 REGF\[6\].RFW.BIT\[24\].FF/Q REGF\[6\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[24] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.INV2\[0\] DEC1.D2.AND5/X VGND VGND VPWR VPWR REGF\[21\].RFW.INV2\[0\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[18\].RFW.BIT\[17\].OBUF1 REGF\[18\].RFW.BIT\[17\].FF/Q REGF\[18\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[17] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.BIT\[30\].OBUF1 REGF\[19\].RFW.BIT\[30\].FF/Q REGF\[19\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[30] sky130_fd_sc_hd__ebufn_2
XREGF\[2\].RFW.BIT\[1\].OBUF2 REGF\[2\].RFW.BIT\[1\].FF/Q REGF\[2\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[1] sky130_fd_sc_hd__ebufn_2
Xfill_46_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_46_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_46_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_62_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_62_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_62_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[23\].RFW.BIT\[7\].OBUF1 REGF\[23\].RFW.BIT\[7\].FF/Q REGF\[23\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[7] sky130_fd_sc_hd__ebufn_2
XDEC2.D0.ABUF\[2\] RW[2] VGND VGND VPWR VPWR DEC2.D0.AND7/C sky130_fd_sc_hd__clkbuf_2
XREGF\[29\].RFW.BIT\[30\].FF REGF\[29\].RFW.CG\[3\]/GCLK DW[30] VGND VGND VPWR VPWR
+ REGF\[29\].RFW.BIT\[30\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[30\].RFW.BIT\[24\].OBUF2 REGF\[30\].RFW.BIT\[24\].FF/Q REGF\[30\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[24] sky130_fd_sc_hd__ebufn_2
XREGF\[30\].RFW.CG\[3\] CLK REGF\[30\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[30\].RFW.CG\[3\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[14\].RFW.BIT\[2\].OBUF2 REGF\[14\].RFW.BIT\[2\].FF/Q REGF\[14\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[2] sky130_fd_sc_hd__ebufn_2
Xfill_21_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[2\].RFW.BIT\[27\].OBUF1 REGF\[2\].RFW.BIT\[27\].FF/Q REGF\[2\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[27] sky130_fd_sc_hd__ebufn_2
Xfill_14_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[28\].RFW.BIT\[20\].OBUF2 REGF\[28\].RFW.BIT\[20\].FF/Q REGF\[28\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[20] sky130_fd_sc_hd__ebufn_2
XREGF\[20\].RFW.BIT\[22\].OBUF1 REGF\[20\].RFW.BIT\[22\].FF/Q REGF\[20\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[22] sky130_fd_sc_hd__ebufn_2
XREGF\[7\].RFW.BIT\[19\].FF REGF\[7\].RFW.CG\[2\]/GCLK DW[19] VGND VGND VPWR VPWR
+ REGF\[7\].RFW.BIT\[19\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[4\].RFW.BIT\[1\].OBUF2 REGF\[4\].RFW.BIT\[1\].FF/Q REGF\[4\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[1] sky130_fd_sc_hd__ebufn_2
Xtap_36_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.BIT\[21\].FF REGF\[3\].RFW.CG\[2\]/GCLK DW[21] VGND VGND VPWR VPWR
+ REGF\[3\].RFW.BIT\[21\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[5\].RFW.BIT\[12\].OBUF1 REGF\[5\].RFW.BIT\[12\].FF/Q REGF\[5\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[12] sky130_fd_sc_hd__ebufn_2
Xfill_16_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_16_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.BIT\[28\].OBUF2 REGF\[6\].RFW.BIT\[28\].FF/Q REGF\[6\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[28] sky130_fd_sc_hd__ebufn_2
XREGF\[25\].RFW.BIT\[7\].OBUF1 REGF\[25\].RFW.BIT\[7\].FF/Q REGF\[25\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[7] sky130_fd_sc_hd__ebufn_2
Xfill_32_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_62_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_32_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_32_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_55_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[16\].RFW.INV2\[1\] DEC1.D2.AND0/Y VGND VGND VPWR VPWR REGF\[16\].RFW.INV2\[1\]/Y
+ sky130_fd_sc_hd__inv_4
Xtap_48_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[24\].RFW.BIT\[19\].FF REGF\[24\].RFW.CG\[2\]/GCLK DW[19] VGND VGND VPWR VPWR
+ REGF\[24\].RFW.BIT\[19\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[24\].RFW.BIT\[23\].OBUF2 REGF\[24\].RFW.BIT\[23\].FF/Q REGF\[24\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[23] sky130_fd_sc_hd__ebufn_2
XREGF\[20\].RFW.BIT\[21\].FF REGF\[20\].RFW.CG\[2\]/GCLK DW[21] VGND VGND VPWR VPWR
+ REGF\[20\].RFW.BIT\[21\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[16\].RFW.BIT\[2\].OBUF2 REGF\[16\].RFW.BIT\[2\].FF/Q REGF\[16\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[2] sky130_fd_sc_hd__ebufn_2
XREGF\[9\].RFW.BIT\[13\].OBUF2 REGF\[9\].RFW.BIT\[13\].FF/Q REGF\[9\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[13] sky130_fd_sc_hd__ebufn_2
Xfill_57_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_57_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_57_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_57_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_57_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_4_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_4_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_57_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[1\].RFW.BIT\[15\].OBUF1 REGF\[1\].RFW.BIT\[15\].FF/Q REGF\[1\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[15] sky130_fd_sc_hd__ebufn_2
XREGF\[14\].RFW.BIT\[21\].OBUF1 REGF\[14\].RFW.BIT\[21\].FF/Q REGF\[14\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[21] sky130_fd_sc_hd__ebufn_2
XREGF\[6\].RFW.BIT\[1\].OBUF2 REGF\[6\].RFW.BIT\[1\].FF/Q REGF\[6\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[1] sky130_fd_sc_hd__ebufn_2
XREGF\[7\].RFW.CG\[3\] CLK REGF\[7\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[7\].RFW.CG\[3\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[19\].RFW.BIT\[26\].FF REGF\[19\].RFW.CG\[3\]/GCLK DW[26] VGND VGND VPWR VPWR
+ REGF\[19\].RFW.BIT\[26\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[31\].RFW.BIT\[31\].FF REGF\[31\].RFW.CG\[3\]/GCLK DW[31] VGND VGND VPWR VPWR
+ REGF\[31\].RFW.BIT\[31\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[20\].RFW.BIT\[26\].OBUF2 REGF\[20\].RFW.BIT\[26\].FF/Q REGF\[20\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[26] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[7\].OBUF1 REGF\[27\].RFW.BIT\[7\].FF/Q REGF\[27\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[7] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[16\].OBUF2 REGF\[5\].RFW.BIT\[16\].FF/Q REGF\[5\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[16] sky130_fd_sc_hd__ebufn_2
XREGF\[12\].RFW.INV1\[2\] DEC0.D1.AND4/X VGND VGND VPWR VPWR REGF\[12\].RFW.INV1\[2\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[18\].RFW.BIT\[22\].OBUF2 REGF\[18\].RFW.BIT\[22\].FF/Q REGF\[18\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[22] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.BIT\[2\].OBUF2 REGF\[18\].RFW.BIT\[2\].FF/Q REGF\[18\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[2] sky130_fd_sc_hd__ebufn_2
XREGF\[10\].RFW.BIT\[24\].OBUF1 REGF\[10\].RFW.BIT\[24\].FF/Q REGF\[10\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[24] sky130_fd_sc_hd__ebufn_2
XREGF\[23\].RFW.BIT\[11\].OBUF2 REGF\[23\].RFW.BIT\[11\].FF/Q REGF\[23\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[11] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.INV1\[3\] DEC0.D3.AND4/X VGND VGND VPWR VPWR REGF\[28\].RFW.INV1\[3\]/Y
+ sky130_fd_sc_hd__inv_4
Xtap_34_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.CG\[0\] CLK REGF\[6\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[6\].RFW.CG\[0\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_27_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[5\].OBUF1 REGF\[20\].RFW.BIT\[5\].FF/Q REGF\[20\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[5] sky130_fd_sc_hd__ebufn_2
XREGF\[8\].RFW.BIT\[1\].OBUF2 REGF\[8\].RFW.BIT\[1\].FF/Q REGF\[8\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[1] sky130_fd_sc_hd__ebufn_2
Xfill_27_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_27_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_27_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_27_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_43_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_43_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_43_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_43_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_43_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[11\].RFW.BIT\[0\].OBUF2 REGF\[11\].RFW.BIT\[0\].FF/Q REGF\[11\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[0] sky130_fd_sc_hd__ebufn_2
XREGF\[1\].RFW.BIT\[19\].OBUF2 REGF\[1\].RFW.BIT\[19\].FF/Q REGF\[1\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[19] sky130_fd_sc_hd__ebufn_2
XREGF\[10\].RFW.BIT\[17\].FF REGF\[10\].RFW.CG\[2\]/GCLK DW[17] VGND VGND VPWR VPWR
+ REGF\[10\].RFW.BIT\[17\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[4\].RFW.BIT\[27\].FF REGF\[4\].RFW.CG\[3\]/GCLK DW[27] VGND VGND VPWR VPWR
+ REGF\[4\].RFW.BIT\[27\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[29\].RFW.BIT\[7\].OBUF1 REGF\[29\].RFW.BIT\[7\].FF/Q REGF\[29\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[7] sky130_fd_sc_hd__ebufn_2
XREGF\[14\].RFW.BIT\[25\].OBUF2 REGF\[14\].RFW.BIT\[25\].FF/Q REGF\[14\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[25] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[11\].FF REGF\[16\].RFW.CG\[1\]/GCLK DW[11] VGND VGND VPWR VPWR
+ REGF\[16\].RFW.BIT\[11\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_55_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_48_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[17\].RFW.BIT\[10\].OBUF2 REGF\[17\].RFW.BIT\[10\].FF/Q REGF\[17\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[10] sky130_fd_sc_hd__ebufn_2
XREGF\[22\].RFW.BIT\[5\].OBUF1 REGF\[22\].RFW.BIT\[5\].FF/Q REGF\[22\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[5] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.BIT\[27\].FF REGF\[21\].RFW.CG\[3\]/GCLK DW[27] VGND VGND VPWR VPWR
+ REGF\[21\].RFW.BIT\[27\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[27\].RFW.BIT\[21\].FF REGF\[27\].RFW.CG\[2\]/GCLK DW[21] VGND VGND VPWR VPWR
+ REGF\[27\].RFW.BIT\[21\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[13\].RFW.BIT\[0\].OBUF2 REGF\[13\].RFW.BIT\[0\].FF/Q REGF\[13\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[0] sky130_fd_sc_hd__ebufn_2
XREGF\[10\].RFW.BIT\[28\].OBUF2 REGF\[10\].RFW.BIT\[28\].FF/Q REGF\[10\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[28] sky130_fd_sc_hd__ebufn_2
Xfill_13_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[9\].OBUF2 REGF\[20\].RFW.BIT\[9\].FF/Q REGF\[20\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[9] sky130_fd_sc_hd__ebufn_2
Xfill_13_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_13_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_13_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[1\].RFW.BIT\[20\].OBUF2 REGF\[1\].RFW.BIT\[20\].FF/Q REGF\[1\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[20] sky130_fd_sc_hd__ebufn_2
Xfill_13_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[13\].RFW.BIT\[13\].OBUF2 REGF\[13\].RFW.BIT\[13\].FF/Q REGF\[13\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[13] sky130_fd_sc_hd__ebufn_2
Xtap_32_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgenblk1.RFW0.INV2\[2\] DEC1.D0.AND0/Y VGND VGND VPWR VPWR genblk1.RFW0.INV2\[2\]/Y
+ sky130_fd_sc_hd__inv_4
Xtap_25_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[1\].RFW.BIT\[12\].FF REGF\[1\].RFW.CG\[1\]/GCLK DW[12] VGND VGND VPWR VPWR
+ REGF\[1\].RFW.BIT\[12\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_18_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_38_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_38_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_38_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.BIT\[27\].OBUF1 REGF\[31\].RFW.BIT\[27\].FF/Q REGF\[31\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[27] sky130_fd_sc_hd__ebufn_2
Xgenblk1.RFW0.BIT\[0\].OBUF1 genblk1.RFW0.TIE\[0\]/LO genblk1.RFW0.INV1\[0\]/Y VGND
+ VGND VPWR VPWR DA[0] sky130_fd_sc_hd__ebufn_2
XDEC1.D0.AND1 DEC1.D0.AND7/C DEC1.D0.AND7/B DEC1.D0.AND7/A DEC1.D0.AND7/D VGND VGND
+ VPWR VPWR DEC1.D0.AND1/X sky130_fd_sc_hd__and4bb_2
Xfill_54_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_54_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_54_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_1_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[24\].RFW.BIT\[5\].OBUF1 REGF\[24\].RFW.BIT\[5\].FF/Q REGF\[24\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[5] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.BIT\[23\].OBUF1 REGF\[29\].RFW.BIT\[23\].FF/Q REGF\[29\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[23] sky130_fd_sc_hd__ebufn_2
XREGF\[15\].RFW.BIT\[0\].OBUF2 REGF\[15\].RFW.BIT\[0\].FF/Q REGF\[15\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[0] sky130_fd_sc_hd__ebufn_2
Xfill_60_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_53_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_46_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[22\].RFW.BIT\[9\].OBUF2 REGF\[22\].RFW.BIT\[9\].FF/Q REGF\[22\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[9] sky130_fd_sc_hd__ebufn_2
Xfill_39_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC0.D1.AND3 DEC0.D1.AND7/C DEC0.D1.AND7/B DEC0.D1.AND7/A DEC0.D1.AND7/D VGND VGND
+ VPWR VPWR DEC0.D1.AND3/X sky130_fd_sc_hd__and4b_2
XREGF\[25\].RFW.BIT\[26\].OBUF1 REGF\[25\].RFW.BIT\[26\].FF/Q REGF\[25\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[26] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.BIT\[17\].FF REGF\[17\].RFW.CG\[2\]/GCLK DW[17] VGND VGND VPWR VPWR
+ REGF\[17\].RFW.BIT\[17\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[30\].RFW.BIT\[15\].OBUF1 REGF\[30\].RFW.BIT\[15\].FF/Q REGF\[30\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[15] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[5\].OBUF1 REGF\[26\].RFW.BIT\[5\].FF/Q REGF\[26\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[5] sky130_fd_sc_hd__ebufn_2
Xtap_4_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_24_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_24_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_24_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XREGF\[28\].RFW.BIT\[11\].OBUF1 REGF\[28\].RFW.BIT\[11\].FF/Q REGF\[28\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[11] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.BIT\[0\].OBUF2 REGF\[17\].RFW.BIT\[0\].FF/Q REGF\[17\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[0] sky130_fd_sc_hd__ebufn_2
Xgenblk1.RFW0.BIT\[4\].OBUF2 genblk1.RFW0.TIE\[4\]/LO genblk1.RFW0.INV2\[0\]/Y VGND
+ VGND VPWR VPWR DB[4] sky130_fd_sc_hd__ebufn_2
Xfill_40_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_40_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_40_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[24\].RFW.BIT\[9\].OBUF2 REGF\[24\].RFW.BIT\[9\].FF/Q REGF\[24\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[9] sky130_fd_sc_hd__ebufn_2
Xfill_49_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_49_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[28\].RFW.BIT\[27\].FF REGF\[28\].RFW.CG\[3\]/GCLK DW[27] VGND VGND VPWR VPWR
+ REGF\[28\].RFW.BIT\[27\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_49_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_49_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_49_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[29\].RFW.BIT\[27\].OBUF2 REGF\[29\].RFW.BIT\[27\].FF/Q REGF\[29\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[27] sky130_fd_sc_hd__ebufn_2
Xfill_49_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[21\].RFW.BIT\[29\].OBUF1 REGF\[21\].RFW.BIT\[29\].FF/Q REGF\[21\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[29] sky130_fd_sc_hd__ebufn_2
Xfill_18_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.BIT\[19\].OBUF1 REGF\[6\].RFW.BIT\[19\].FF/Q REGF\[6\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[19] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.BIT\[25\].OBUF1 REGF\[19\].RFW.BIT\[25\].FF/Q REGF\[19\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[25] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.BIT\[5\].OBUF1 REGF\[28\].RFW.BIT\[5\].FF/Q REGF\[28\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[5] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[14\].OBUF1 REGF\[24\].RFW.BIT\[14\].FF/Q REGF\[24\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[14] sky130_fd_sc_hd__ebufn_2
XREGF\[2\].RFW.BIT\[18\].FF REGF\[2\].RFW.CG\[2\]/GCLK DW[18] VGND VGND VPWR VPWR
+ REGF\[2\].RFW.BIT\[18\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_51_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_44_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[8\].RFW.BIT\[12\].FF REGF\[8\].RFW.CG\[1\]/GCLK DW[12] VGND VGND VPWR VPWR
+ REGF\[8\].RFW.BIT\[12\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_37_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[19\].RFW.BIT\[0\].OBUF2 REGF\[19\].RFW.BIT\[0\].FF/Q REGF\[19\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[0] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[9\].OBUF2 REGF\[26\].RFW.BIT\[9\].FF/Q REGF\[26\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[9] sky130_fd_sc_hd__ebufn_2
XREGF\[30\].RFW.BIT\[19\].OBUF2 REGF\[30\].RFW.BIT\[19\].FF/Q REGF\[30\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[19] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.BIT\[3\].OBUF1 REGF\[21\].RFW.BIT\[3\].FF/Q REGF\[21\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[3] sky130_fd_sc_hd__ebufn_2
Xfill_10_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_10_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[15\].RFW.BIT\[28\].OBUF1 REGF\[15\].RFW.BIT\[28\].FF/Q REGF\[15\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[28] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.BIT\[15\].OBUF2 REGF\[28\].RFW.BIT\[15\].FF/Q REGF\[28\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[15] sky130_fd_sc_hd__ebufn_2
Xfill_19_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_19_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_19_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_19_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_19_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[17\].OBUF1 REGF\[20\].RFW.BIT\[17\].FF/Q REGF\[20\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[17] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.BIT\[30\].OBUF1 REGF\[21\].RFW.BIT\[30\].FF/Q REGF\[21\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[30] sky130_fd_sc_hd__ebufn_2
Xtap_2_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[25\].RFW.BIT\[12\].FF REGF\[25\].RFW.CG\[1\]/GCLK DW[12] VGND VGND VPWR VPWR
+ REGF\[25\].RFW.BIT\[12\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_35_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_35_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_35_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_35_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.BIT\[20\].OBUF1 REGF\[6\].RFW.BIT\[20\].FF/Q REGF\[6\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[20] sky130_fd_sc_hd__ebufn_2
Xfill_51_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_51_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_51_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.BIT\[13\].OBUF1 REGF\[18\].RFW.BIT\[13\].FF/Q REGF\[18\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[13] sky130_fd_sc_hd__ebufn_2
Xfill_51_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_51_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_7_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_7_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_7_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_7_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[14\].RFW.BIT\[25\].FF REGF\[14\].RFW.CG\[3\]/GCLK DW[25] VGND VGND VPWR VPWR
+ REGF\[14\].RFW.BIT\[25\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[30\].RFW.BIT\[28\].FF REGF\[30\].RFW.CG\[3\]/GCLK DW[28] VGND VGND VPWR VPWR
+ REGF\[30\].RFW.BIT\[28\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[19\].RFW.BIT\[29\].OBUF2 REGF\[19\].RFW.BIT\[29\].FF/Q REGF\[19\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[29] sky130_fd_sc_hd__ebufn_2
Xfill_30_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[28\].RFW.BIT\[9\].OBUF2 REGF\[28\].RFW.BIT\[9\].FF/Q REGF\[28\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[9] sky130_fd_sc_hd__ebufn_2
Xfill_23_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[23\].RFW.BIT\[3\].OBUF1 REGF\[23\].RFW.BIT\[3\].FF/Q REGF\[23\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[3] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[18\].OBUF2 REGF\[24\].RFW.BIT\[18\].FF/Q REGF\[24\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[18] sky130_fd_sc_hd__ebufn_2
Xfill_16_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[25\].RFW.BIT\[31\].OBUF2 REGF\[25\].RFW.BIT\[31\].FF/Q REGF\[25\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[31] sky130_fd_sc_hd__ebufn_2
XREGF\[30\].RFW.BIT\[20\].OBUF2 REGF\[30\].RFW.BIT\[20\].FF/Q REGF\[30\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[20] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.BIT\[1\].FF REGF\[17\].RFW.CG\[0\]/GCLK DW[1] VGND VGND VPWR VPWR
+ REGF\[17\].RFW.BIT\[1\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[4\].RFW.INV2\[3\] DEC1.D0.AND4/X VGND VGND VPWR VPWR REGF\[4\].RFW.INV2\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[2\].RFW.BIT\[23\].OBUF1 REGF\[2\].RFW.BIT\[23\].FF/Q REGF\[2\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[23] sky130_fd_sc_hd__ebufn_2
XREGF\[14\].RFW.BIT\[16\].OBUF1 REGF\[14\].RFW.BIT\[16\].FF/Q REGF\[14\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[16] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.BIT\[7\].OBUF2 REGF\[21\].RFW.BIT\[7\].FF/Q REGF\[21\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[7] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[3\].FF REGF\[16\].RFW.CG\[0\]/GCLK DW[3] VGND VGND VPWR VPWR
+ REGF\[16\].RFW.BIT\[3\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[24\].RFW.INV2\[1\] DEC1.D3.AND0/Y VGND VGND VPWR VPWR REGF\[24\].RFW.INV2\[1\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_21_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_21_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.BIT\[24\].OBUF2 REGF\[6\].RFW.BIT\[24\].FF/Q REGF\[6\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[24] sky130_fd_sc_hd__ebufn_2
XREGF\[15\].RFW.BIT\[5\].FF REGF\[15\].RFW.CG\[0\]/GCLK DW[5] VGND VGND VPWR VPWR
+ REGF\[15\].RFW.BIT\[5\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[25\].RFW.BIT\[3\].OBUF1 REGF\[25\].RFW.BIT\[3\].FF/Q REGF\[25\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[3] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.BIT\[17\].OBUF2 REGF\[18\].RFW.BIT\[17\].FF/Q REGF\[18\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[17] sky130_fd_sc_hd__ebufn_2
XREGF\[9\].RFW.BIT\[18\].FF REGF\[9\].RFW.CG\[2\]/GCLK DW[18] VGND VGND VPWR VPWR
+ REGF\[9\].RFW.BIT\[18\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[19\].RFW.BIT\[30\].OBUF2 REGF\[19\].RFW.BIT\[30\].FF/Q REGF\[19\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[30] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[20\].FF REGF\[5\].RFW.CG\[2\]/GCLK DW[20] VGND VGND VPWR VPWR
+ REGF\[5\].RFW.BIT\[20\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[11\].RFW.BIT\[10\].FF REGF\[11\].RFW.CG\[1\]/GCLK DW[10] VGND VGND VPWR VPWR
+ REGF\[11\].RFW.BIT\[10\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_0_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_46_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_46_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_46_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[10\].RFW.BIT\[19\].OBUF1 REGF\[10\].RFW.BIT\[19\].FF/Q REGF\[10\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[19] sky130_fd_sc_hd__ebufn_2
Xfill_62_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_62_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_62_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.CG\[2\] CLK REGF\[3\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[3\].RFW.CG\[2\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[14\].RFW.BIT\[7\].FF REGF\[14\].RFW.CG\[0\]/GCLK DW[7] VGND VGND VPWR VPWR
+ REGF\[14\].RFW.BIT\[7\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[1\].RFW.BIT\[11\].OBUF1 REGF\[1\].RFW.BIT\[11\].FF/Q REGF\[1\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[11] sky130_fd_sc_hd__ebufn_2
XREGF\[23\].RFW.BIT\[7\].OBUF2 REGF\[23\].RFW.BIT\[7\].FF/Q REGF\[23\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[7] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[18\].FF REGF\[26\].RFW.CG\[2\]/GCLK DW[18] VGND VGND VPWR VPWR
+ REGF\[26\].RFW.BIT\[18\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[29\].RFW.BIT\[3\].FF REGF\[29\].RFW.CG\[0\]/GCLK DW[3] VGND VGND VPWR VPWR
+ REGF\[29\].RFW.BIT\[3\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_21_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[2\].RFW.BIT\[27\].OBUF2 REGF\[2\].RFW.BIT\[27\].FF/Q REGF\[2\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[27] sky130_fd_sc_hd__ebufn_2
XREGF\[20\].RFW.INV1\[2\] DEC0.D2.AND4/X VGND VGND VPWR VPWR REGF\[20\].RFW.INV1\[2\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[22\].RFW.BIT\[20\].FF REGF\[22\].RFW.CG\[2\]/GCLK DW[20] VGND VGND VPWR VPWR
+ REGF\[22\].RFW.BIT\[20\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[13\].RFW.BIT\[9\].FF REGF\[13\].RFW.CG\[1\]/GCLK DW[9] VGND VGND VPWR VPWR
+ REGF\[13\].RFW.BIT\[9\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[29\].RFW.CG\[1\] CLK REGF\[29\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[29\].RFW.CG\[1\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[20\].RFW.BIT\[22\].OBUF2 REGF\[20\].RFW.BIT\[22\].FF/Q REGF\[20\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[22] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[3\].OBUF1 REGF\[27\].RFW.BIT\[3\].FF/Q REGF\[27\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[3] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.BIT\[5\].FF REGF\[28\].RFW.CG\[0\]/GCLK DW[5] VGND VGND VPWR VPWR
+ REGF\[28\].RFW.BIT\[5\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[5\].RFW.BIT\[12\].OBUF2 REGF\[5\].RFW.BIT\[12\].FF/Q REGF\[5\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[12] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.INV2\[2\] DEC1.D2.AND3/X VGND VGND VPWR VPWR REGF\[19\].RFW.INV2\[2\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[10\].RFW.BIT\[20\].OBUF1 REGF\[10\].RFW.BIT\[20\].FF/Q REGF\[10\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[20] sky130_fd_sc_hd__ebufn_2
Xfill_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_16_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[25\].RFW.BIT\[7\].OBUF2 REGF\[25\].RFW.BIT\[7\].FF/Q REGF\[25\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[7] sky130_fd_sc_hd__ebufn_2
XREGF\[20\].RFW.BIT\[1\].OBUF1 REGF\[20\].RFW.BIT\[1\].FF/Q REGF\[20\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[1] sky130_fd_sc_hd__ebufn_2
Xfill_32_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[27\].RFW.BIT\[7\].FF REGF\[27\].RFW.CG\[0\]/GCLK DW[7] VGND VGND VPWR VPWR
+ REGF\[27\].RFW.BIT\[7\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_62_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_32_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_32_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_55_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_48_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_57_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_57_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_57_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_57_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_4_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_4_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_57_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_57_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[26\].RFW.BIT\[9\].FF REGF\[26\].RFW.CG\[1\]/GCLK DW[9] VGND VGND VPWR VPWR
+ REGF\[26\].RFW.BIT\[9\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[1\].RFW.BIT\[15\].OBUF2 REGF\[1\].RFW.BIT\[15\].FF/Q REGF\[1\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[15] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.BIT\[3\].OBUF1 REGF\[29\].RFW.BIT\[3\].FF/Q REGF\[29\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[3] sky130_fd_sc_hd__ebufn_2
XREGF\[14\].RFW.BIT\[21\].OBUF2 REGF\[14\].RFW.BIT\[21\].FF/Q REGF\[14\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[21] sky130_fd_sc_hd__ebufn_2
XREGF\[15\].RFW.INV1\[3\] DEC0.D1.AND7/X VGND VGND VPWR VPWR REGF\[15\].RFW.INV1\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[17\].RFW.CG\[1\] CLK REGF\[17\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[17\].RFW.CG\[1\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[29\].RFW.BIT\[18\].OBUF1 REGF\[29\].RFW.BIT\[18\].FF/Q REGF\[29\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[18] sky130_fd_sc_hd__ebufn_2
XREGF\[6\].RFW.BIT\[26\].FF REGF\[6\].RFW.CG\[3\]/GCLK DW[26] VGND VGND VPWR VPWR
+ REGF\[6\].RFW.BIT\[26\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[12\].RFW.BIT\[16\].FF REGF\[12\].RFW.CG\[2\]/GCLK DW[16] VGND VGND VPWR VPWR
+ REGF\[12\].RFW.BIT\[16\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[27\].RFW.BIT\[7\].OBUF2 REGF\[27\].RFW.BIT\[7\].FF/Q REGF\[27\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[7] sky130_fd_sc_hd__ebufn_2
XREGF\[22\].RFW.BIT\[1\].OBUF1 REGF\[22\].RFW.BIT\[1\].FF/Q REGF\[22\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[1] sky130_fd_sc_hd__ebufn_2
Xfill_12_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.BIT\[10\].FF REGF\[18\].RFW.CG\[1\]/GCLK DW[10] VGND VGND VPWR VPWR
+ REGF\[18\].RFW.BIT\[10\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[10\].RFW.BIT\[24\].OBUF2 REGF\[10\].RFW.BIT\[24\].FF/Q REGF\[10\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[24] sky130_fd_sc_hd__ebufn_2
Xtap_34_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[5\].OBUF2 REGF\[20\].RFW.BIT\[5\].FF/Q REGF\[20\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[5] sky130_fd_sc_hd__ebufn_2
Xfill_27_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_27_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_27_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[23\].RFW.BIT\[26\].FF REGF\[23\].RFW.CG\[3\]/GCLK DW[26] VGND VGND VPWR VPWR
+ REGF\[23\].RFW.BIT\[26\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_27_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_27_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_43_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[29\].RFW.BIT\[20\].FF REGF\[29\].RFW.CG\[2\]/GCLK DW[20] VGND VGND VPWR VPWR
+ REGF\[29\].RFW.BIT\[20\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_43_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_43_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_43_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_43_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.BIT\[23\].OBUF1 REGF\[31\].RFW.BIT\[23\].FF/Q REGF\[31\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[23] sky130_fd_sc_hd__ebufn_2
Xtap_60_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[29\].RFW.BIT\[7\].OBUF2 REGF\[29\].RFW.BIT\[7\].FF/Q REGF\[29\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[7] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[1\].OBUF1 REGF\[24\].RFW.BIT\[1\].FF/Q REGF\[24\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[1] sky130_fd_sc_hd__ebufn_2
Xfill_48_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.INV2\[0\] DEC1.D0.AND6/X VGND VGND VPWR VPWR REGF\[6\].RFW.INV2\[0\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_3_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.BIT\[11\].FF REGF\[3\].RFW.CG\[1\]/GCLK DW[11] VGND VGND VPWR VPWR
+ REGF\[3\].RFW.BIT\[11\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[22\].RFW.BIT\[5\].OBUF2 REGF\[22\].RFW.BIT\[5\].FF/Q REGF\[22\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[5] sky130_fd_sc_hd__ebufn_2
XREGF\[7\].RFW.BIT\[27\].OBUF1 REGF\[7\].RFW.BIT\[27\].FF/Q REGF\[7\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[27] sky130_fd_sc_hd__ebufn_2
Xfill_5_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[25\].RFW.BIT\[22\].OBUF1 REGF\[25\].RFW.BIT\[22\].FF/Q REGF\[25\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[22] sky130_fd_sc_hd__ebufn_2
XREGF\[20\].RFW.BIT\[11\].FF REGF\[20\].RFW.CG\[1\]/GCLK DW[11] VGND VGND VPWR VPWR
+ REGF\[20\].RFW.BIT\[11\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_13_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[26\].RFW.BIT\[1\].OBUF1 REGF\[26\].RFW.BIT\[1\].FF/Q REGF\[26\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[1] sky130_fd_sc_hd__ebufn_2
XREGF\[30\].RFW.BIT\[11\].OBUF1 REGF\[30\].RFW.BIT\[11\].FF/Q REGF\[30\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[11] sky130_fd_sc_hd__ebufn_2
Xfill_13_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_13_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_13_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_38_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[2\].RFW.INV1\[1\] DEC0.D0.AND2/X VGND VGND VPWR VPWR REGF\[2\].RFW.INV1\[1\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_38_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_38_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.BIT\[27\].OBUF2 REGF\[31\].RFW.BIT\[27\].FF/Q REGF\[31\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[27] sky130_fd_sc_hd__ebufn_2
XDEC1.D0.AND2 DEC1.D0.AND7/C DEC1.D0.AND7/A DEC1.D0.AND7/B DEC1.D0.AND7/D VGND VGND
+ VPWR VPWR DEC1.D0.AND2/X sky130_fd_sc_hd__and4bb_2
Xgenblk1.RFW0.BIT\[0\].OBUF2 genblk1.RFW0.TIE\[4\]/LO genblk1.RFW0.INV2\[0\]/Y VGND
+ VGND VPWR VPWR DB[0] sky130_fd_sc_hd__ebufn_2
Xfill_54_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_54_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[19\].RFW.BIT\[16\].FF REGF\[19\].RFW.CG\[2\]/GCLK DW[16] VGND VGND VPWR VPWR
+ REGF\[19\].RFW.BIT\[16\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_54_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[24\].RFW.BIT\[5\].OBUF2 REGF\[24\].RFW.BIT\[5\].FF/Q REGF\[24\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[5] sky130_fd_sc_hd__ebufn_2
XREGF\[31\].RFW.BIT\[21\].FF REGF\[31\].RFW.CG\[2\]/GCLK DW[21] VGND VGND VPWR VPWR
+ REGF\[31\].RFW.BIT\[21\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[29\].RFW.BIT\[23\].OBUF2 REGF\[29\].RFW.BIT\[23\].FF/Q REGF\[29\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[23] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.BIT\[25\].OBUF1 REGF\[21\].RFW.BIT\[25\].FF/Q REGF\[21\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[25] sky130_fd_sc_hd__ebufn_2
Xfill_60_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.BIT\[15\].OBUF1 REGF\[6\].RFW.BIT\[15\].FF/Q REGF\[6\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[15] sky130_fd_sc_hd__ebufn_2
Xfill_53_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[11\].RFW.BIT\[0\].FF REGF\[11\].RFW.CG\[0\]/GCLK DW[0] VGND VGND VPWR VPWR
+ REGF\[11\].RFW.BIT\[0\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[19\].RFW.BIT\[21\].OBUF1 REGF\[19\].RFW.BIT\[21\].FF/Q REGF\[19\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[21] sky130_fd_sc_hd__ebufn_2
Xfill_46_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_39_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[28\].RFW.BIT\[1\].OBUF1 REGF\[28\].RFW.BIT\[1\].FF/Q REGF\[28\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[1] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[10\].OBUF1 REGF\[24\].RFW.BIT\[10\].FF/Q REGF\[24\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[10] sky130_fd_sc_hd__ebufn_2
Xfill_1_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC0.D1.AND4 DEC0.D1.AND7/A DEC0.D1.AND7/B DEC0.D1.AND7/C DEC0.D1.AND7/D VGND VGND
+ VPWR VPWR DEC0.D1.AND4/X sky130_fd_sc_hd__and4bb_2
XREGF\[10\].RFW.BIT\[2\].FF REGF\[10\].RFW.CG\[0\]/GCLK DW[2] VGND VGND VPWR VPWR
+ REGF\[10\].RFW.BIT\[2\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[25\].RFW.BIT\[26\].OBUF2 REGF\[25\].RFW.BIT\[26\].FF/Q REGF\[25\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[26] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[5\].OBUF2 REGF\[26\].RFW.BIT\[5\].FF/Q REGF\[26\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[5] sky130_fd_sc_hd__ebufn_2
XREGF\[30\].RFW.BIT\[15\].OBUF2 REGF\[30\].RFW.BIT\[15\].FF/Q REGF\[30\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[15] sky130_fd_sc_hd__ebufn_2
Xtap_4_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[2\].RFW.BIT\[18\].OBUF1 REGF\[2\].RFW.BIT\[18\].FF/Q REGF\[2\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[18] sky130_fd_sc_hd__ebufn_2
XREGF\[3\].RFW.BIT\[31\].OBUF1 REGF\[3\].RFW.BIT\[31\].FF/Q REGF\[3\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[31] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.BIT\[17\].FF REGF\[4\].RFW.CG\[2\]/GCLK DW[17] VGND VGND VPWR VPWR
+ REGF\[4\].RFW.BIT\[17\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_24_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[15\].RFW.BIT\[24\].OBUF1 REGF\[15\].RFW.BIT\[24\].FF/Q REGF\[15\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[24] sky130_fd_sc_hd__ebufn_2
Xfill_24_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[28\].RFW.BIT\[11\].OBUF2 REGF\[28\].RFW.BIT\[11\].FF/Q REGF\[28\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[11] sky130_fd_sc_hd__ebufn_2
XREGF\[20\].RFW.BIT\[13\].OBUF1 REGF\[20\].RFW.BIT\[13\].FF/Q REGF\[20\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[13] sky130_fd_sc_hd__ebufn_2
Xfill_40_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_40_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_40_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_49_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_49_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_49_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_49_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_49_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[24\].RFW.BIT\[0\].FF REGF\[24\].RFW.CG\[0\]/GCLK DW[0] VGND VGND VPWR VPWR
+ REGF\[24\].RFW.BIT\[0\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[21\].RFW.BIT\[29\].OBUF2 REGF\[21\].RFW.BIT\[29\].FF/Q REGF\[21\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[29] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.BIT\[17\].FF REGF\[21\].RFW.CG\[2\]/GCLK DW[17] VGND VGND VPWR VPWR
+ REGF\[21\].RFW.BIT\[17\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[6\].RFW.BIT\[19\].OBUF2 REGF\[6\].RFW.BIT\[19\].FF/Q REGF\[6\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[19] sky130_fd_sc_hd__ebufn_2
XDEC2.TIE VGND VGND VPWR VPWR DEC2.TIE/HI DEC2.TIE/LO sky130_fd_sc_hd__conb_1
XREGF\[17\].RFW.INV1\[0\] DEC0.D2.AND1/X VGND VGND VPWR VPWR REGF\[17\].RFW.INV1\[0\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[19\].RFW.BIT\[25\].OBUF2 REGF\[19\].RFW.BIT\[25\].FF/Q REGF\[19\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[25] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[11\].FF REGF\[27\].RFW.CG\[1\]/GCLK DW[11] VGND VGND VPWR VPWR
+ REGF\[27\].RFW.BIT\[11\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[23\].RFW.BIT\[2\].FF REGF\[23\].RFW.CG\[0\]/GCLK DW[2] VGND VGND VPWR VPWR
+ REGF\[23\].RFW.BIT\[2\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[28\].RFW.BIT\[5\].OBUF2 REGF\[28\].RFW.BIT\[5\].FF/Q REGF\[28\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[5] sky130_fd_sc_hd__ebufn_2
XREGF\[11\].RFW.BIT\[27\].OBUF1 REGF\[11\].RFW.BIT\[27\].FF/Q REGF\[11\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[27] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[14\].OBUF2 REGF\[24\].RFW.BIT\[14\].FF/Q REGF\[24\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[14] sky130_fd_sc_hd__ebufn_2
Xfill_51_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_44_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[30\].RFW.BIT\[8\].OBUF1 REGF\[30\].RFW.BIT\[8\].FF/Q REGF\[30\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[8] sky130_fd_sc_hd__ebufn_2
Xfill_37_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[16\].RFW.BIT\[24\].FF REGF\[16\].RFW.CG\[3\]/GCLK DW[24] VGND VGND VPWR VPWR
+ REGF\[16\].RFW.BIT\[24\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[14\].RFW.BIT\[12\].OBUF1 REGF\[14\].RFW.BIT\[12\].FF/Q REGF\[14\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[12] sky130_fd_sc_hd__ebufn_2
XREGF\[22\].RFW.BIT\[4\].FF REGF\[22\].RFW.CG\[0\]/GCLK DW[4] VGND VGND VPWR VPWR
+ REGF\[22\].RFW.BIT\[4\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[21\].RFW.BIT\[3\].OBUF2 REGF\[21\].RFW.BIT\[3\].FF/Q REGF\[21\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[3] sky130_fd_sc_hd__ebufn_2
Xfill_10_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_10_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[15\].RFW.BIT\[28\].OBUF2 REGF\[15\].RFW.BIT\[28\].FF/Q REGF\[15\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[28] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.CG\[3\] CLK REGF\[26\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[26\].RFW.CG\[3\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_19_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_19_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_19_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_19_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[21\].RFW.BIT\[6\].FF REGF\[21\].RFW.CG\[0\]/GCLK DW[6] VGND VGND VPWR VPWR
+ REGF\[21\].RFW.BIT\[6\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_19_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[17\].OBUF2 REGF\[20\].RFW.BIT\[17\].FF/Q REGF\[20\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[17] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.BIT\[30\].OBUF2 REGF\[21\].RFW.BIT\[30\].FF/Q REGF\[21\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[30] sky130_fd_sc_hd__ebufn_2
Xtap_2_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_35_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[6\].RFW.BIT\[20\].OBUF2 REGF\[6\].RFW.BIT\[20\].FF/Q REGF\[6\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[20] sky130_fd_sc_hd__ebufn_2
Xfill_51_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_51_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[18\].RFW.BIT\[13\].OBUF2 REGF\[18\].RFW.BIT\[13\].FF/Q REGF\[18\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[13] sky130_fd_sc_hd__ebufn_2
Xfill_51_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_51_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[7\].RFW.BIT\[1\].FF REGF\[7\].RFW.CG\[0\]/GCLK DW[1] VGND VGND VPWR VPWR REGF\[7\].RFW.BIT\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xfill_51_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[10\].RFW.BIT\[15\].OBUF1 REGF\[10\].RFW.BIT\[15\].FF/Q REGF\[10\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[15] sky130_fd_sc_hd__ebufn_2
Xfill_7_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[8\].FF REGF\[20\].RFW.CG\[1\]/GCLK DW[8] VGND VGND VPWR VPWR
+ REGF\[20\].RFW.BIT\[8\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_7_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_7_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_30_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[25\].RFW.CG\[0\] CLK REGF\[25\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[25\].RFW.CG\[0\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_23_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[23\].RFW.BIT\[3\].OBUF2 REGF\[23\].RFW.BIT\[3\].FF/Q REGF\[23\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[3] sky130_fd_sc_hd__ebufn_2
XREGF\[6\].RFW.BIT\[3\].FF REGF\[6\].RFW.CG\[0\]/GCLK DW[3] VGND VGND VPWR VPWR REGF\[6\].RFW.BIT\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[1\].RFW.BIT\[25\].FF REGF\[1\].RFW.CG\[3\]/GCLK DW[25] VGND VGND VPWR VPWR
+ REGF\[1\].RFW.BIT\[25\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_16_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[11\].RFW.INV2\[1\] DEC1.D1.AND3/X VGND VGND VPWR VPWR REGF\[11\].RFW.INV2\[1\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[2\].RFW.BIT\[23\].OBUF2 REGF\[2\].RFW.BIT\[23\].FF/Q REGF\[2\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[23] sky130_fd_sc_hd__ebufn_2
XREGF\[14\].RFW.BIT\[16\].OBUF2 REGF\[14\].RFW.BIT\[16\].FF/Q REGF\[14\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[16] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.INV2\[2\] DEC1.D3.AND3/X VGND VGND VPWR VPWR REGF\[27\].RFW.INV2\[2\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[5\].RFW.BIT\[5\].FF REGF\[5\].RFW.CG\[0\]/GCLK DW[5] VGND VGND VPWR VPWR REGF\[5\].RFW.BIT\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xfill_42_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[28\].RFW.BIT\[17\].FF REGF\[28\].RFW.CG\[2\]/GCLK DW[17] VGND VGND VPWR VPWR
+ REGF\[28\].RFW.BIT\[17\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[14\].RFW.CG\[3\] CLK REGF\[14\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[14\].RFW.CG\[3\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[4\].RFW.BIT\[7\].FF REGF\[4\].RFW.CG\[0\]/GCLK DW[7] VGND VGND VPWR VPWR REGF\[4\].RFW.BIT\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xfill_21_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xtap_4_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[25\].RFW.BIT\[3\].OBUF2 REGF\[25\].RFW.BIT\[3\].FF/Q REGF\[25\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[3] sky130_fd_sc_hd__ebufn_2
Xtap_0_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_46_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_46_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_46_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[10\].RFW.BIT\[19\].OBUF2 REGF\[10\].RFW.BIT\[19\].FF/Q REGF\[10\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[19] sky130_fd_sc_hd__ebufn_2
Xfill_62_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[3\].RFW.BIT\[9\].FF REGF\[3\].RFW.CG\[1\]/GCLK DW[9] VGND VGND VPWR VPWR REGF\[3\].RFW.BIT\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xfill_62_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_62_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[23\].RFW.INV1\[3\] DEC0.D2.AND7/X VGND VGND VPWR VPWR REGF\[23\].RFW.INV1\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[13\].RFW.CG\[0\] CLK REGF\[13\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[13\].RFW.CG\[0\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[1\].RFW.BIT\[11\].OBUF2 REGF\[1\].RFW.BIT\[11\].FF/Q REGF\[1\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[11] sky130_fd_sc_hd__ebufn_2
Xfill_11_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[26\].RFW.BIT\[29\].OBUF1 REGF\[26\].RFW.BIT\[29\].FF/Q REGF\[26\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[29] sky130_fd_sc_hd__ebufn_2
XREGF\[31\].RFW.BIT\[18\].OBUF1 REGF\[31\].RFW.BIT\[18\].FF/Q REGF\[31\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[18] sky130_fd_sc_hd__ebufn_2
Xfill_21_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_14_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[29\].RFW.BIT\[14\].OBUF1 REGF\[29\].RFW.BIT\[14\].FF/Q REGF\[29\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[14] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[3\].OBUF2 REGF\[27\].RFW.BIT\[3\].FF/Q REGF\[27\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[3] sky130_fd_sc_hd__ebufn_2
XREGF\[10\].RFW.BIT\[20\].OBUF2 REGF\[10\].RFW.BIT\[20\].FF/Q REGF\[10\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[20] sky130_fd_sc_hd__ebufn_2
Xfill_16_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XDEC2.D2.ABUF\[1\] RW[1] VGND VGND VPWR VPWR DEC2.D2.AND7/B sky130_fd_sc_hd__clkbuf_2
XREGF\[8\].RFW.BIT\[25\].FF REGF\[8\].RFW.CG\[3\]/GCLK DW[25] VGND VGND VPWR VPWR
+ REGF\[8\].RFW.BIT\[25\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[14\].RFW.BIT\[15\].FF REGF\[14\].RFW.CG\[1\]/GCLK DW[15] VGND VGND VPWR VPWR
+ REGF\[14\].RFW.BIT\[15\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[20\].RFW.BIT\[1\].OBUF2 REGF\[20\].RFW.BIT\[1\].FF/Q REGF\[20\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[1] sky130_fd_sc_hd__ebufn_2
Xtap_62_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_32_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_32_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_32_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[30\].RFW.BIT\[18\].FF REGF\[30\].RFW.CG\[2\]/GCLK DW[18] VGND VGND VPWR VPWR
+ REGF\[30\].RFW.BIT\[18\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_55_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_48_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[25\].RFW.BIT\[17\].OBUF1 REGF\[25\].RFW.BIT\[17\].FF/Q REGF\[25\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[17] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[30\].OBUF1 REGF\[26\].RFW.BIT\[30\].FF/Q REGF\[26\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[30] sky130_fd_sc_hd__ebufn_2
Xfill_57_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_57_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_57_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_57_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_4_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDEC1.D3.AND0 DEC1.D3.AND7/A DEC1.D3.AND7/B DEC1.D3.AND7/C DEC1.D3.AND7/D VGND VGND
+ VPWR VPWR DEC1.D3.AND0/Y sky130_fd_sc_hd__nor4b_2
Xfill_57_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[29\].RFW.BIT\[3\].OBUF2 REGF\[29\].RFW.BIT\[3\].FF/Q REGF\[29\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[3] sky130_fd_sc_hd__ebufn_2
XREGF\[25\].RFW.BIT\[25\].FF REGF\[25\].RFW.CG\[3\]/GCLK DW[25] VGND VGND VPWR VPWR
+ REGF\[25\].RFW.BIT\[25\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[31\].RFW.BIT\[6\].OBUF1 REGF\[31\].RFW.BIT\[6\].FF/Q REGF\[31\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[6] sky130_fd_sc_hd__ebufn_2
Xgenblk1.RFW0.TIE\[5\] VGND VGND VPWR VPWR genblk1.RFW0.TIE\[5\]/HI genblk1.RFW0.TIE\[5\]/LO
+ sky130_fd_sc_hd__conb_1
XREGF\[29\].RFW.BIT\[18\].OBUF2 REGF\[29\].RFW.BIT\[18\].FF/Q REGF\[29\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[18] sky130_fd_sc_hd__ebufn_2
XREGF\[22\].RFW.BIT\[1\].OBUF2 REGF\[22\].RFW.BIT\[1\].FF/Q REGF\[22\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[1] sky130_fd_sc_hd__ebufn_2
Xfill_12_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[7\].RFW.BIT\[23\].OBUF1 REGF\[7\].RFW.BIT\[23\].FF/Q REGF\[7\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[23] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.BIT\[16\].OBUF1 REGF\[19\].RFW.BIT\[16\].FF/Q REGF\[19\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[16] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[10\].FF REGF\[5\].RFW.CG\[1\]/GCLK DW[10] VGND VGND VPWR VPWR
+ REGF\[5\].RFW.BIT\[10\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_34_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_27_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_27_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_27_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_27_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_27_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_43_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_43_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_43_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_43_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_43_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xtap_60_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.BIT\[23\].OBUF2 REGF\[31\].RFW.BIT\[23\].FF/Q REGF\[31\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[23] sky130_fd_sc_hd__ebufn_2
Xtap_53_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[9\].RFW.INV2\[1\] DEC1.D1.AND1/X VGND VGND VPWR VPWR REGF\[9\].RFW.INV2\[1\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[22\].RFW.BIT\[10\].FF REGF\[22\].RFW.CG\[1\]/GCLK DW[10] VGND VGND VPWR VPWR
+ REGF\[22\].RFW.BIT\[10\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[24\].RFW.BIT\[1\].OBUF2 REGF\[24\].RFW.BIT\[1\].FF/Q REGF\[24\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[1] sky130_fd_sc_hd__ebufn_2
XREGF\[3\].RFW.BIT\[26\].OBUF1 REGF\[3\].RFW.BIT\[26\].FF/Q REGF\[3\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[26] sky130_fd_sc_hd__ebufn_2
XREGF\[15\].RFW.BIT\[19\].OBUF1 REGF\[15\].RFW.BIT\[19\].FF/Q REGF\[15\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[19] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.BIT\[21\].OBUF1 REGF\[21\].RFW.BIT\[21\].FF/Q REGF\[21\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[21] sky130_fd_sc_hd__ebufn_2
XREGF\[6\].RFW.BIT\[11\].OBUF1 REGF\[6\].RFW.BIT\[11\].FF/Q REGF\[6\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[11] sky130_fd_sc_hd__ebufn_2
XREGF\[11\].RFW.BIT\[23\].FF REGF\[11\].RFW.CG\[2\]/GCLK DW[23] VGND VGND VPWR VPWR
+ REGF\[11\].RFW.BIT\[23\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[7\].RFW.BIT\[27\].OBUF2 REGF\[7\].RFW.BIT\[27\].FF/Q REGF\[7\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[27] sky130_fd_sc_hd__ebufn_2
Xfill_5_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_5_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_8_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[25\].RFW.BIT\[22\].OBUF2 REGF\[25\].RFW.BIT\[22\].FF/Q REGF\[25\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[22] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.INV1\[2\] DEC0.D0.AND5/X VGND VGND VPWR VPWR REGF\[5\].RFW.INV1\[2\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[26\].RFW.BIT\[1\].OBUF2 REGF\[26\].RFW.BIT\[1\].FF/Q REGF\[26\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[1] sky130_fd_sc_hd__ebufn_2
XREGF\[30\].RFW.BIT\[11\].OBUF2 REGF\[30\].RFW.BIT\[11\].FF/Q REGF\[30\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[11] sky130_fd_sc_hd__ebufn_2
Xfill_13_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_13_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_13_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[2\].RFW.BIT\[14\].OBUF1 REGF\[2\].RFW.BIT\[14\].FF/Q REGF\[2\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[14] sky130_fd_sc_hd__ebufn_2
XDEC1.D3.ABUF\[2\] RB[2] VGND VGND VPWR VPWR DEC1.D3.AND7/C sky130_fd_sc_hd__clkbuf_2
Xtap_32_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[15\].RFW.BIT\[20\].OBUF1 REGF\[15\].RFW.BIT\[20\].FF/Q REGF\[15\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[20] sky130_fd_sc_hd__ebufn_2
Xtap_25_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_38_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_38_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_38_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC1.D0.AND3 DEC1.D0.AND7/C DEC1.D0.AND7/B DEC1.D0.AND7/A DEC1.D0.AND7/D VGND VGND
+ VPWR VPWR DEC1.D0.AND3/X sky130_fd_sc_hd__and4b_2
XREGF\[1\].RFW.BIT\[0\].FF REGF\[1\].RFW.CG\[0\]/GCLK DW[0] VGND VGND VPWR VPWR REGF\[1\].RFW.BIT\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[30\].RFW.BIT\[1\].FF REGF\[30\].RFW.CG\[0\]/GCLK DW[1] VGND VGND VPWR VPWR
+ REGF\[30\].RFW.BIT\[1\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_54_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_54_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[25\].RFW.INV1\[0\] DEC0.D3.AND1/X VGND VGND VPWR VPWR REGF\[25\].RFW.INV1\[0\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_54_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_1_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.BIT\[16\].FF REGF\[6\].RFW.CG\[2\]/GCLK DW[16] VGND VGND VPWR VPWR
+ REGF\[6\].RFW.BIT\[16\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[21\].RFW.BIT\[25\].OBUF2 REGF\[21\].RFW.BIT\[25\].FF/Q REGF\[21\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[25] sky130_fd_sc_hd__ebufn_2
Xfill_60_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.BIT\[15\].OBUF2 REGF\[6\].RFW.BIT\[15\].FF/Q REGF\[6\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[15] sky130_fd_sc_hd__ebufn_2
Xfill_53_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[19\].RFW.BIT\[21\].OBUF2 REGF\[19\].RFW.BIT\[21\].FF/Q REGF\[19\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[21] sky130_fd_sc_hd__ebufn_2
Xfill_46_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_39_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[28\].RFW.BIT\[1\].OBUF2 REGF\[28\].RFW.BIT\[1\].FF/Q REGF\[28\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[1] sky130_fd_sc_hd__ebufn_2
XREGF\[11\].RFW.BIT\[23\].OBUF1 REGF\[11\].RFW.BIT\[23\].FF/Q REGF\[11\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[23] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[10\].OBUF2 REGF\[24\].RFW.BIT\[10\].FF/Q REGF\[24\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[10] sky130_fd_sc_hd__ebufn_2
Xfill_1_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[30\].RFW.BIT\[4\].OBUF1 REGF\[30\].RFW.BIT\[4\].FF/Q REGF\[30\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[4] sky130_fd_sc_hd__ebufn_2
XREGF\[23\].RFW.BIT\[16\].FF REGF\[23\].RFW.CG\[2\]/GCLK DW[16] VGND VGND VPWR VPWR
+ REGF\[23\].RFW.BIT\[16\].FF/Q sky130_fd_sc_hd__dfxtp_1
XDEC0.D1.AND5 DEC0.D1.AND7/B DEC0.D1.AND7/A DEC0.D1.AND7/C DEC0.D1.AND7/D VGND VGND
+ VPWR VPWR DEC0.D1.AND5/X sky130_fd_sc_hd__and4b_2
XREGF\[22\].RFW.CG\[2\] CLK REGF\[22\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[22\].RFW.CG\[2\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[29\].RFW.BIT\[10\].FF REGF\[29\].RFW.CG\[1\]/GCLK DW[10] VGND VGND VPWR VPWR
+ REGF\[29\].RFW.BIT\[10\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_4_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[2\].RFW.BIT\[18\].OBUF2 REGF\[2\].RFW.BIT\[18\].FF/Q REGF\[2\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[18] sky130_fd_sc_hd__ebufn_2
XREGF\[3\].RFW.BIT\[31\].OBUF2 REGF\[3\].RFW.BIT\[31\].FF/Q REGF\[3\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[31] sky130_fd_sc_hd__ebufn_2
Xfill_24_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.BIT\[29\].FF REGF\[12\].RFW.CG\[3\]/GCLK DW[29] VGND VGND VPWR VPWR
+ REGF\[12\].RFW.BIT\[29\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[15\].RFW.BIT\[24\].OBUF2 REGF\[15\].RFW.BIT\[24\].FF/Q REGF\[15\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[24] sky130_fd_sc_hd__ebufn_2
Xfill_24_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[13\].OBUF2 REGF\[20\].RFW.BIT\[13\].FF/Q REGF\[20\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[13] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.BIT\[23\].FF REGF\[18\].RFW.CG\[2\]/GCLK DW[23] VGND VGND VPWR VPWR
+ REGF\[18\].RFW.BIT\[23\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_40_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_40_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_40_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_30_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_49_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xtap_23_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_49_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_49_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_49_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xtap_16_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_49_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[10\].RFW.BIT\[11\].OBUF1 REGF\[10\].RFW.BIT\[11\].FF/Q REGF\[10\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[11] sky130_fd_sc_hd__ebufn_2
XREGF\[11\].RFW.BIT\[27\].OBUF2 REGF\[11\].RFW.BIT\[27\].FF/Q REGF\[11\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[27] sky130_fd_sc_hd__ebufn_2
Xfill_51_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_44_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[30\].RFW.BIT\[8\].OBUF2 REGF\[30\].RFW.BIT\[8\].FF/Q REGF\[30\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[8] sky130_fd_sc_hd__ebufn_2
Xfill_37_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[14\].RFW.BIT\[12\].OBUF2 REGF\[14\].RFW.BIT\[12\].FF/Q REGF\[14\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[12] sky130_fd_sc_hd__ebufn_2
XREGF\[10\].RFW.CG\[2\] CLK REGF\[10\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[10\].RFW.CG\[2\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[3\].RFW.BIT\[24\].FF REGF\[3\].RFW.CG\[3\]/GCLK DW[24] VGND VGND VPWR VPWR
+ REGF\[3\].RFW.BIT\[24\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_10_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.BIT\[11\].FF REGF\[31\].RFW.CG\[1\]/GCLK DW[11] VGND VGND VPWR VPWR
+ REGF\[31\].RFW.BIT\[11\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_19_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_19_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_19_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_19_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_35_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_35_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.INV1\[3\] DEC0.D3.AND7/X VGND VGND VPWR VPWR REGF\[31\].RFW.INV1\[3\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_51_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_51_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_51_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_51_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_51_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[10\].RFW.BIT\[15\].OBUF2 REGF\[10\].RFW.BIT\[15\].FF/Q REGF\[10\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[15] sky130_fd_sc_hd__ebufn_2
XREGF\[20\].RFW.BIT\[24\].FF REGF\[20\].RFW.CG\[3\]/GCLK DW[24] VGND VGND VPWR VPWR
+ REGF\[20\].RFW.BIT\[24\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_7_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_7_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[14\].RFW.INV2\[2\] DEC1.D1.AND6/X VGND VGND VPWR VPWR REGF\[14\].RFW.INV2\[2\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_23_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_16_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[26\].RFW.BIT\[25\].OBUF1 REGF\[26\].RFW.BIT\[25\].FF/Q REGF\[26\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[25] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.BIT\[29\].FF REGF\[19\].RFW.CG\[3\]/GCLK DW[29] VGND VGND VPWR VPWR
+ REGF\[19\].RFW.BIT\[29\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[31\].RFW.BIT\[14\].OBUF1 REGF\[31\].RFW.BIT\[14\].FF/Q REGF\[31\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[14] sky130_fd_sc_hd__ebufn_2
XREGF\[15\].RFW.BIT\[31\].FF REGF\[15\].RFW.CG\[3\]/GCLK DW[31] VGND VGND VPWR VPWR
+ REGF\[15\].RFW.BIT\[31\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[29\].RFW.BIT\[10\].OBUF1 REGF\[29\].RFW.BIT\[10\].FF/Q REGF\[29\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[10] sky130_fd_sc_hd__ebufn_2
Xfill_42_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_35_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xtap_4_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[22\].RFW.BIT\[28\].OBUF1 REGF\[22\].RFW.BIT\[28\].FF/Q REGF\[22\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[28] sky130_fd_sc_hd__ebufn_2
XREGF\[10\].RFW.INV1\[3\] DEC0.D1.AND2/X VGND VGND VPWR VPWR REGF\[10\].RFW.INV1\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[7\].RFW.BIT\[18\].OBUF1 REGF\[7\].RFW.BIT\[18\].FF/Q REGF\[7\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[18] sky130_fd_sc_hd__ebufn_2
XREGF\[8\].RFW.BIT\[31\].OBUF1 REGF\[8\].RFW.BIT\[31\].FF/Q REGF\[8\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[31] sky130_fd_sc_hd__ebufn_2
Xfill_46_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_46_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_46_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_62_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[25\].RFW.BIT\[13\].OBUF1 REGF\[25\].RFW.BIT\[13\].FF/Q REGF\[25\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[13] sky130_fd_sc_hd__ebufn_2
Xfill_62_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_62_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_11_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_11_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[16\].RFW.BIT\[14\].FF REGF\[16\].RFW.CG\[1\]/GCLK DW[14] VGND VGND VPWR VPWR
+ REGF\[16\].RFW.BIT\[14\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[26\].RFW.BIT\[29\].OBUF2 REGF\[26\].RFW.BIT\[29\].FF/Q REGF\[26\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[29] sky130_fd_sc_hd__ebufn_2
XREGF\[31\].RFW.BIT\[18\].OBUF2 REGF\[31\].RFW.BIT\[18\].FF/Q REGF\[31\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[18] sky130_fd_sc_hd__ebufn_2
XREGF\[31\].RFW.BIT\[2\].OBUF1 REGF\[31\].RFW.BIT\[2\].FF/Q REGF\[31\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[2] sky130_fd_sc_hd__ebufn_2
Xfill_21_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_14_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[16\].RFW.BIT\[27\].OBUF1 REGF\[16\].RFW.BIT\[27\].FF/Q REGF\[16\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[27] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.BIT\[14\].OBUF2 REGF\[29\].RFW.BIT\[14\].FF/Q REGF\[29\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[14] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.BIT\[16\].OBUF1 REGF\[21\].RFW.BIT\[16\].FF/Q REGF\[21\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[16] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[24\].FF REGF\[27\].RFW.CG\[3\]/GCLK DW[24] VGND VGND VPWR VPWR
+ REGF\[27\].RFW.BIT\[24\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[19\].RFW.BIT\[12\].OBUF1 REGF\[19\].RFW.BIT\[12\].FF/Q REGF\[19\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[12] sky130_fd_sc_hd__ebufn_2
XREGF\[1\].RFW.INV2\[0\] DEC1.D0.AND1/X VGND VGND VPWR VPWR REGF\[1\].RFW.INV2\[0\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_16_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_16_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xtap_62_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_32_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_32_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_32_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_48_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[25\].RFW.BIT\[17\].OBUF2 REGF\[25\].RFW.BIT\[17\].FF/Q REGF\[25\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[17] sky130_fd_sc_hd__ebufn_2
XREGF\[1\].RFW.BIT\[15\].FF REGF\[1\].RFW.CG\[1\]/GCLK DW[15] VGND VGND VPWR VPWR
+ REGF\[1\].RFW.BIT\[15\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[26\].RFW.BIT\[30\].OBUF2 REGF\[26\].RFW.BIT\[30\].FF/Q REGF\[26\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[30] sky130_fd_sc_hd__ebufn_2
Xfill_57_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_57_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_57_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_4_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC1.D3.AND1 DEC1.D3.AND7/C DEC1.D3.AND7/B DEC1.D3.AND7/A DEC1.D3.AND7/D VGND VGND
+ VPWR VPWR DEC1.D3.AND1/X sky130_fd_sc_hd__and4bb_2
Xfill_57_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_57_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[3\].RFW.BIT\[22\].OBUF1 REGF\[3\].RFW.BIT\[22\].FF/Q REGF\[3\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[22] sky130_fd_sc_hd__ebufn_2
XREGF\[15\].RFW.BIT\[15\].OBUF1 REGF\[15\].RFW.BIT\[15\].FF/Q REGF\[15\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[15] sky130_fd_sc_hd__ebufn_2
XREGF\[31\].RFW.BIT\[6\].OBUF2 REGF\[31\].RFW.BIT\[6\].FF/Q REGF\[31\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[6] sky130_fd_sc_hd__ebufn_2
XDEC2.D0.ABUF\[0\] RW[0] VGND VGND VPWR VPWR DEC2.D0.AND7/A sky130_fd_sc_hd__clkbuf_2
XREGF\[30\].RFW.CG\[1\] CLK REGF\[30\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[30\].RFW.CG\[1\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_12_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XREGF\[7\].RFW.BIT\[23\].OBUF2 REGF\[7\].RFW.BIT\[23\].FF/Q REGF\[7\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[23] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.BIT\[16\].OBUF2 REGF\[19\].RFW.BIT\[16\].FF/Q REGF\[19\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[16] sky130_fd_sc_hd__ebufn_2
XREGF\[12\].RFW.BIT\[31\].OBUF1 REGF\[12\].RFW.BIT\[31\].FF/Q REGF\[12\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[31] sky130_fd_sc_hd__ebufn_2
XREGF\[11\].RFW.BIT\[18\].OBUF1 REGF\[11\].RFW.BIT\[18\].FF/Q REGF\[11\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[18] sky130_fd_sc_hd__ebufn_2
Xtap_34_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[13\].RFW.BIT\[22\].FF REGF\[13\].RFW.CG\[2\]/GCLK DW[22] VGND VGND VPWR VPWR
+ REGF\[13\].RFW.BIT\[22\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_27_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_27_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_27_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_27_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[2\].RFW.BIT\[10\].OBUF1 REGF\[2\].RFW.BIT\[10\].FF/Q REGF\[2\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[10] sky130_fd_sc_hd__ebufn_2
Xfill_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_43_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_43_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_43_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_43_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_60_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_53_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_46_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.BIT\[26\].OBUF2 REGF\[3\].RFW.BIT\[26\].FF/Q REGF\[3\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[26] sky130_fd_sc_hd__ebufn_2
XREGF\[15\].RFW.BIT\[19\].OBUF2 REGF\[15\].RFW.BIT\[19\].FF/Q REGF\[15\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[19] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.BIT\[21\].OBUF2 REGF\[21\].RFW.BIT\[21\].FF/Q REGF\[21\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[21] sky130_fd_sc_hd__ebufn_2
Xfill_17_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[6\].RFW.BIT\[11\].OBUF2 REGF\[6\].RFW.BIT\[11\].FF/Q REGF\[6\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[11] sky130_fd_sc_hd__ebufn_2
XREGF\[7\].RFW.CG\[1\] CLK REGF\[7\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[7\].RFW.CG\[1\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[8\].RFW.INV1\[3\] DEC0.D1.AND0/Y VGND VGND VPWR VPWR REGF\[8\].RFW.INV1\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[8\].RFW.BIT\[15\].FF REGF\[8\].RFW.CG\[1\]/GCLK DW[15] VGND VGND VPWR VPWR
+ REGF\[8\].RFW.BIT\[15\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_5_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfill_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_5_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[30\].RFW.BIT\[0\].OBUF1 REGF\[30\].RFW.BIT\[0\].FF/Q REGF\[30\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[0] sky130_fd_sc_hd__ebufn_2
Xfill_8_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[12\].RFW.INV1\[0\] DEC0.D1.AND4/X VGND VGND VPWR VPWR REGF\[12\].RFW.INV1\[0\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_13_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_13_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[28\].RFW.INV1\[1\] DEC0.D3.AND4/X VGND VGND VPWR VPWR REGF\[28\].RFW.INV1\[1\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[2\].RFW.BIT\[14\].OBUF2 REGF\[2\].RFW.BIT\[14\].FF/Q REGF\[2\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[14] sky130_fd_sc_hd__ebufn_2
Xtap_32_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_25_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[15\].RFW.BIT\[20\].OBUF2 REGF\[15\].RFW.BIT\[20\].FF/Q REGF\[15\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[20] sky130_fd_sc_hd__ebufn_2
Xtap_18_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[19\].RFW.BIT\[0\].FF REGF\[19\].RFW.CG\[0\]/GCLK DW[0] VGND VGND VPWR VPWR
+ REGF\[19\].RFW.BIT\[0\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[25\].RFW.BIT\[15\].FF REGF\[25\].RFW.CG\[1\]/GCLK DW[15] VGND VGND VPWR VPWR
+ REGF\[25\].RFW.BIT\[15\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_38_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_38_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_38_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDEC1.D0.AND4 DEC1.D0.AND7/A DEC1.D0.AND7/B DEC1.D0.AND7/C DEC1.D0.AND7/D VGND VGND
+ VPWR VPWR DEC1.D0.AND4/X sky130_fd_sc_hd__and4bb_2
Xfill_54_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_54_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_54_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.BIT\[2\].FF REGF\[18\].RFW.CG\[0\]/GCLK DW[2] VGND VGND VPWR VPWR
+ REGF\[18\].RFW.BIT\[2\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[14\].RFW.BIT\[28\].FF REGF\[14\].RFW.CG\[3\]/GCLK DW[28] VGND VGND VPWR VPWR
+ REGF\[14\].RFW.BIT\[28\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[10\].RFW.BIT\[30\].FF REGF\[10\].RFW.CG\[3\]/GCLK DW[30] VGND VGND VPWR VPWR
+ REGF\[10\].RFW.BIT\[30\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_53_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_46_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC1.D1.ABUF\[1\] RB[1] VGND VGND VPWR VPWR DEC1.D1.AND7/B sky130_fd_sc_hd__clkbuf_2
XREGF\[11\].RFW.BIT\[23\].OBUF2 REGF\[11\].RFW.BIT\[23\].FF/Q REGF\[11\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[23] sky130_fd_sc_hd__ebufn_2
Xfill_1_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[17\].RFW.BIT\[4\].FF REGF\[17\].RFW.CG\[0\]/GCLK DW[4] VGND VGND VPWR VPWR
+ REGF\[17\].RFW.BIT\[4\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[30\].RFW.BIT\[4\].OBUF2 REGF\[30\].RFW.BIT\[4\].FF/Q REGF\[30\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[4] sky130_fd_sc_hd__ebufn_2
XDEC0.D1.AND6 DEC0.D1.AND7/A DEC0.D1.AND7/B DEC0.D1.AND7/C DEC0.D1.AND7/D VGND VGND
+ VPWR VPWR DEC0.D1.AND6/X sky130_fd_sc_hd__and4b_2
XREGF\[16\].RFW.BIT\[6\].FF REGF\[16\].RFW.CG\[0\]/GCLK DW[6] VGND VGND VPWR VPWR
+ REGF\[16\].RFW.BIT\[6\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_24_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_24_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_40_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_40_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_40_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[15\].RFW.BIT\[8\].FF REGF\[15\].RFW.CG\[1\]/GCLK DW[8] VGND VGND VPWR VPWR
+ REGF\[15\].RFW.BIT\[8\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[22\].RFW.INV2\[2\] DEC1.D2.AND6/X VGND VGND VPWR VPWR REGF\[22\].RFW.INV2\[2\]/Y
+ sky130_fd_sc_hd__inv_4
Xtap_30_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_49_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_49_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_49_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_49_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgenblk1.RFW0.INV2\[0\] DEC1.D0.AND0/Y VGND VGND VPWR VPWR genblk1.RFW0.INV2\[0\]/Y
+ sky130_fd_sc_hd__inv_4
Xtap_16_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_49_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[5\].RFW.BIT\[23\].FF REGF\[5\].RFW.CG\[2\]/GCLK DW[23] VGND VGND VPWR VPWR
+ REGF\[5\].RFW.BIT\[23\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[11\].RFW.BIT\[13\].FF REGF\[11\].RFW.CG\[1\]/GCLK DW[13] VGND VGND VPWR VPWR
+ REGF\[11\].RFW.BIT\[13\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_9_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[10\].RFW.BIT\[11\].OBUF2 REGF\[10\].RFW.BIT\[11\].FF/Q REGF\[10\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[11] sky130_fd_sc_hd__ebufn_2
XREGF\[8\].RFW.BIT\[26\].OBUF1 REGF\[8\].RFW.BIT\[26\].FF/Q REGF\[8\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[26] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[21\].OBUF1 REGF\[26\].RFW.BIT\[21\].FF/Q REGF\[26\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[21] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.BIT\[6\].FF REGF\[29\].RFW.CG\[0\]/GCLK DW[6] VGND VGND VPWR VPWR
+ REGF\[29\].RFW.BIT\[6\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_51_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_44_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[31\].RFW.BIT\[10\].OBUF1 REGF\[31\].RFW.BIT\[10\].FF/Q REGF\[31\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[10] sky130_fd_sc_hd__ebufn_2
XREGF\[22\].RFW.BIT\[23\].FF REGF\[22\].RFW.CG\[2\]/GCLK DW[23] VGND VGND VPWR VPWR
+ REGF\[22\].RFW.BIT\[23\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_37_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_2_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[28\].RFW.BIT\[8\].FF REGF\[28\].RFW.CG\[1\]/GCLK DW[8] VGND VGND VPWR VPWR
+ REGF\[28\].RFW.BIT\[8\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_10_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[4\].RFW.BIT\[29\].OBUF1 REGF\[4\].RFW.BIT\[29\].FF/Q REGF\[4\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[29] sky130_fd_sc_hd__ebufn_2
Xfill_19_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_19_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_19_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[17\].RFW.BIT\[30\].FF REGF\[17\].RFW.CG\[3\]/GCLK DW[30] VGND VGND VPWR VPWR
+ REGF\[17\].RFW.BIT\[30\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_2_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[22\].RFW.BIT\[24\].OBUF1 REGF\[22\].RFW.BIT\[24\].FF/Q REGF\[22\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[24] sky130_fd_sc_hd__ebufn_2
Xfill_35_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_35_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[7\].RFW.BIT\[14\].OBUF1 REGF\[7\].RFW.BIT\[14\].FF/Q REGF\[7\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[14] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.INV2\[3\] DEC1.D2.AND1/X VGND VGND VPWR VPWR REGF\[17\].RFW.INV2\[3\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_51_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_51_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_51_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_51_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_51_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_7_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_16_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[26\].RFW.BIT\[25\].OBUF2 REGF\[26\].RFW.BIT\[25\].FF/Q REGF\[26\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[25] sky130_fd_sc_hd__ebufn_2
Xfill_25_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC0.D2.ABUF\[2\] RA[2] VGND VGND VPWR VPWR DEC0.D2.AND7/C sky130_fd_sc_hd__clkbuf_2
XREGF\[31\].RFW.BIT\[14\].OBUF2 REGF\[31\].RFW.BIT\[14\].FF/Q REGF\[31\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[14] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.BIT\[30\].OBUF1 REGF\[4\].RFW.BIT\[30\].FF/Q REGF\[4\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[30] sky130_fd_sc_hd__ebufn_2
XREGF\[3\].RFW.BIT\[17\].OBUF1 REGF\[3\].RFW.BIT\[17\].FF/Q REGF\[3\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[17] sky130_fd_sc_hd__ebufn_2
XREGF\[6\].RFW.BIT\[29\].FF REGF\[6\].RFW.CG\[3\]/GCLK DW[29] VGND VGND VPWR VPWR
+ REGF\[6\].RFW.BIT\[29\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[12\].RFW.BIT\[19\].FF REGF\[12\].RFW.CG\[2\]/GCLK DW[19] VGND VGND VPWR VPWR
+ REGF\[12\].RFW.BIT\[19\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[16\].RFW.BIT\[23\].OBUF1 REGF\[16\].RFW.BIT\[23\].FF/Q REGF\[16\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[23] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.BIT\[10\].OBUF2 REGF\[29\].RFW.BIT\[10\].FF/Q REGF\[29\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[10] sky130_fd_sc_hd__ebufn_2
XREGF\[2\].RFW.BIT\[31\].FF REGF\[2\].RFW.CG\[3\]/GCLK DW[31] VGND VGND VPWR VPWR
+ REGF\[2\].RFW.BIT\[31\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_42_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[21\].RFW.BIT\[12\].OBUF1 REGF\[21\].RFW.BIT\[12\].FF/Q REGF\[21\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[12] sky130_fd_sc_hd__ebufn_2
Xfill_35_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[18\].RFW.BIT\[13\].FF REGF\[18\].RFW.CG\[1\]/GCLK DW[13] VGND VGND VPWR VPWR
+ REGF\[18\].RFW.BIT\[13\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_28_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_21_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_4_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[22\].RFW.BIT\[28\].OBUF2 REGF\[22\].RFW.BIT\[28\].FF/Q REGF\[22\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[28] sky130_fd_sc_hd__ebufn_2
XREGF\[7\].RFW.BIT\[18\].OBUF2 REGF\[7\].RFW.BIT\[18\].FF/Q REGF\[7\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[18] sky130_fd_sc_hd__ebufn_2
XREGF\[8\].RFW.BIT\[31\].OBUF2 REGF\[8\].RFW.BIT\[31\].FF/Q REGF\[8\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[31] sky130_fd_sc_hd__ebufn_2
XREGF\[23\].RFW.BIT\[29\].FF REGF\[23\].RFW.CG\[3\]/GCLK DW[29] VGND VGND VPWR VPWR
+ REGF\[23\].RFW.BIT\[29\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_46_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_46_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xtap_0_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_46_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[29\].RFW.BIT\[23\].FF REGF\[29\].RFW.CG\[2\]/GCLK DW[23] VGND VGND VPWR VPWR
+ REGF\[29\].RFW.BIT\[23\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[12\].RFW.BIT\[26\].OBUF1 REGF\[12\].RFW.BIT\[26\].FF/Q REGF\[12\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[26] sky130_fd_sc_hd__ebufn_2
XREGF\[25\].RFW.BIT\[13\].OBUF2 REGF\[25\].RFW.BIT\[13\].FF/Q REGF\[25\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[13] sky130_fd_sc_hd__ebufn_2
Xfill_62_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_62_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_62_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_11_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_11_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[15\].RFW.BIT\[11\].OBUF1 REGF\[15\].RFW.BIT\[11\].FF/Q REGF\[15\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[11] sky130_fd_sc_hd__ebufn_2
XREGF\[31\].RFW.BIT\[2\].OBUF2 REGF\[31\].RFW.BIT\[2\].FF/Q REGF\[31\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[2] sky130_fd_sc_hd__ebufn_2
XREGF\[3\].RFW.BIT\[14\].FF REGF\[3\].RFW.CG\[1\]/GCLK DW[14] VGND VGND VPWR VPWR
+ REGF\[3\].RFW.BIT\[14\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_21_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgenblk1.RFW0.BIT\[27\].OBUF1 genblk1.RFW0.TIE\[3\]/LO genblk1.RFW0.INV1\[3\]/Y VGND
+ VGND VPWR VPWR DA[27] sky130_fd_sc_hd__ebufn_2
Xfill_14_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC2.D2.AND0 DEC2.D2.AND7/A DEC2.D2.AND7/B DEC2.D2.AND7/C DEC2.D2.AND7/D VGND VGND
+ VPWR VPWR DEC2.D2.AND0/Y sky130_fd_sc_hd__nor4b_2
XREGF\[16\].RFW.BIT\[27\].OBUF2 REGF\[16\].RFW.BIT\[27\].FF/Q REGF\[16\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[27] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.BIT\[16\].OBUF2 REGF\[21\].RFW.BIT\[16\].FF/Q REGF\[21\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[16] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.INV2\[1\] DEC1.D0.AND4/X VGND VGND VPWR VPWR REGF\[4\].RFW.INV2\[1\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[19\].RFW.BIT\[12\].OBUF2 REGF\[19\].RFW.BIT\[12\].FF/Q REGF\[19\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[12] sky130_fd_sc_hd__ebufn_2
Xfill_16_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[14\].FF REGF\[20\].RFW.CG\[1\]/GCLK DW[14] VGND VGND VPWR VPWR
+ REGF\[20\].RFW.BIT\[14\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[4\].RFW.CG\[3\] CLK REGF\[4\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[4\].RFW.CG\[3\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[11\].RFW.BIT\[14\].OBUF1 REGF\[11\].RFW.BIT\[14\].FF/Q REGF\[11\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[14] sky130_fd_sc_hd__ebufn_2
Xfill_16_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_32_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_32_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_32_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_62_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_48_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_57_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_57_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_57_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC1.D3.AND2 DEC1.D3.AND7/C DEC1.D3.AND7/A DEC1.D3.AND7/B DEC1.D3.AND7/D VGND VGND
+ VPWR VPWR DEC1.D3.AND2/X sky130_fd_sc_hd__and4bb_2
Xfill_57_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_57_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[19\].RFW.BIT\[19\].FF REGF\[19\].RFW.CG\[2\]/GCLK DW[19] VGND VGND VPWR VPWR
+ REGF\[19\].RFW.BIT\[19\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[9\].RFW.BIT\[31\].FF REGF\[9\].RFW.CG\[3\]/GCLK DW[31] VGND VGND VPWR VPWR
+ REGF\[9\].RFW.BIT\[31\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[15\].RFW.BIT\[21\].FF REGF\[15\].RFW.CG\[2\]/GCLK DW[21] VGND VGND VPWR VPWR
+ REGF\[15\].RFW.BIT\[21\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[12\].RFW.BIT\[1\].FF REGF\[12\].RFW.CG\[0\]/GCLK DW[1] VGND VGND VPWR VPWR
+ REGF\[12\].RFW.BIT\[1\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[3\].RFW.BIT\[22\].OBUF2 REGF\[3\].RFW.BIT\[22\].FF/Q REGF\[3\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[22] sky130_fd_sc_hd__ebufn_2
XREGF\[31\].RFW.BIT\[24\].FF REGF\[31\].RFW.CG\[3\]/GCLK DW[24] VGND VGND VPWR VPWR
+ REGF\[31\].RFW.BIT\[24\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[15\].RFW.BIT\[15\].OBUF2 REGF\[15\].RFW.BIT\[15\].FF/Q REGF\[15\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[15] sky130_fd_sc_hd__ebufn_2
XREGF\[3\].RFW.CG\[0\] CLK REGF\[3\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[3\].RFW.CG\[0\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[11\].RFW.BIT\[3\].FF REGF\[11\].RFW.CG\[0\]/GCLK DW[3] VGND VGND VPWR VPWR
+ REGF\[11\].RFW.BIT\[3\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[20\].RFW.INV1\[0\] DEC0.D2.AND4/X VGND VGND VPWR VPWR REGF\[20\].RFW.INV1\[0\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[26\].RFW.BIT\[31\].FF REGF\[26\].RFW.CG\[3\]/GCLK DW[31] VGND VGND VPWR VPWR
+ REGF\[26\].RFW.BIT\[31\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_12_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[10\].RFW.BIT\[5\].FF REGF\[10\].RFW.CG\[0\]/GCLK DW[5] VGND VGND VPWR VPWR
+ REGF\[10\].RFW.BIT\[5\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[11\].RFW.BIT\[18\].OBUF2 REGF\[11\].RFW.BIT\[18\].FF/Q REGF\[11\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[18] sky130_fd_sc_hd__ebufn_2
XREGF\[12\].RFW.BIT\[31\].OBUF2 REGF\[12\].RFW.BIT\[31\].FF/Q REGF\[12\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[31] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.INV2\[0\] DEC1.D2.AND3/X VGND VGND VPWR VPWR REGF\[19\].RFW.INV2\[0\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_27_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_27_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_27_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[25\].RFW.BIT\[1\].FF REGF\[25\].RFW.CG\[0\]/GCLK DW[1] VGND VGND VPWR VPWR
+ REGF\[25\].RFW.BIT\[1\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[2\].RFW.BIT\[10\].OBUF2 REGF\[2\].RFW.BIT\[10\].FF/Q REGF\[2\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[10] sky130_fd_sc_hd__ebufn_2
Xfill_43_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_43_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[27\].RFW.BIT\[28\].OBUF1 REGF\[27\].RFW.BIT\[28\].FF/Q REGF\[27\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[28] sky130_fd_sc_hd__ebufn_2
Xfill_43_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_60_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_53_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.CG\[2\] CLK REGF\[18\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[18\].RFW.CG\[2\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_46_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_39_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[24\].RFW.BIT\[3\].FF REGF\[24\].RFW.CG\[0\]/GCLK DW[3] VGND VGND VPWR VPWR
+ REGF\[24\].RFW.BIT\[3\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_17_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_17_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XREGF\[27\].RFW.BIT\[14\].FF REGF\[27\].RFW.CG\[1\]/GCLK DW[14] VGND VGND VPWR VPWR
+ REGF\[27\].RFW.BIT\[14\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_33_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[23\].RFW.BIT\[5\].FF REGF\[23\].RFW.CG\[0\]/GCLK DW[5] VGND VGND VPWR VPWR
+ REGF\[23\].RFW.BIT\[5\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[15\].RFW.INV1\[1\] DEC0.D1.AND7/X VGND VGND VPWR VPWR REGF\[15\].RFW.INV1\[1\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_5_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_5_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_5_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[30\].RFW.BIT\[0\].OBUF2 REGF\[30\].RFW.BIT\[0\].FF/Q REGF\[30\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[0] sky130_fd_sc_hd__ebufn_2
XREGF\[9\].RFW.BIT\[0\].FF REGF\[9\].RFW.CG\[0\]/GCLK DW[0] VGND VGND VPWR VPWR REGF\[9\].RFW.BIT\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[16\].RFW.BIT\[27\].FF REGF\[16\].RFW.CG\[3\]/GCLK DW[27] VGND VGND VPWR VPWR
+ REGF\[16\].RFW.BIT\[27\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[22\].RFW.BIT\[7\].FF REGF\[22\].RFW.CG\[0\]/GCLK DW[7] VGND VGND VPWR VPWR
+ REGF\[22\].RFW.BIT\[7\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_10_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_8_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[26\].RFW.BIT\[16\].OBUF1 REGF\[26\].RFW.BIT\[16\].FF/Q REGF\[26\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[16] sky130_fd_sc_hd__ebufn_2
Xfill_13_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[30\].RFW.INV2\[2\] DEC1.D3.AND6/X VGND VGND VPWR VPWR REGF\[30\].RFW.INV2\[2\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[8\].RFW.BIT\[2\].FF REGF\[8\].RFW.CG\[0\]/GCLK DW[2] VGND VGND VPWR VPWR REGF\[8\].RFW.BIT\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xtap_32_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[21\].RFW.BIT\[9\].FF REGF\[21\].RFW.CG\[1\]/GCLK DW[9] VGND VGND VPWR VPWR
+ REGF\[21\].RFW.BIT\[9\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_18_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_38_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_38_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_38_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDEC1.D0.AND5 DEC1.D0.AND7/B DEC1.D0.AND7/A DEC1.D0.AND7/C DEC1.D0.AND7/D VGND VGND
+ VPWR VPWR DEC1.D0.AND5/X sky130_fd_sc_hd__and4b_2
Xfill_54_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_54_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_54_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[7\].RFW.BIT\[4\].FF REGF\[7\].RFW.CG\[0\]/GCLK DW[4] VGND VGND VPWR VPWR REGF\[7\].RFW.BIT\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[22\].RFW.BIT\[19\].OBUF1 REGF\[22\].RFW.BIT\[19\].FF/Q REGF\[22\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[19] sky130_fd_sc_hd__ebufn_2
XREGF\[8\].RFW.BIT\[22\].OBUF1 REGF\[8\].RFW.BIT\[22\].FF/Q REGF\[8\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[22] sky130_fd_sc_hd__ebufn_2
Xfill_46_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.BIT\[6\].FF REGF\[6\].RFW.CG\[0\]/GCLK DW[6] VGND VGND VPWR VPWR REGF\[6\].RFW.BIT\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[1\].RFW.BIT\[28\].FF REGF\[1\].RFW.CG\[3\]/GCLK DW[28] VGND VGND VPWR VPWR
+ REGF\[1\].RFW.BIT\[28\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_1_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[7\].RFW.BIT\[22\].FF REGF\[7\].RFW.CG\[2\]/GCLK DW[22] VGND VGND VPWR VPWR
+ REGF\[7\].RFW.BIT\[22\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[13\].RFW.BIT\[12\].FF REGF\[13\].RFW.CG\[1\]/GCLK DW[12] VGND VGND VPWR VPWR
+ REGF\[13\].RFW.BIT\[12\].FF/Q sky130_fd_sc_hd__dfxtp_1
XDEC0.D1.AND7 DEC0.D1.AND7/A DEC0.D1.AND7/B DEC0.D1.AND7/C DEC0.D1.AND7/D VGND VGND
+ VPWR VPWR DEC0.D1.AND7/X sky130_fd_sc_hd__and4_2
XREGF\[5\].RFW.BIT\[8\].FF REGF\[5\].RFW.CG\[1\]/GCLK DW[8] VGND VGND VPWR VPWR REGF\[5\].RFW.BIT\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xfill_58_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[25\].RFW.INV2\[3\] DEC1.D3.AND1/X VGND VGND VPWR VPWR REGF\[25\].RFW.INV2\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[4\].RFW.BIT\[25\].OBUF1 REGF\[4\].RFW.BIT\[25\].FF/Q REGF\[4\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[25] sky130_fd_sc_hd__ebufn_2
Xfill_24_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[24\].RFW.BIT\[22\].FF REGF\[24\].RFW.CG\[2\]/GCLK DW[22] VGND VGND VPWR VPWR
+ REGF\[24\].RFW.BIT\[22\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[16\].RFW.BIT\[18\].OBUF1 REGF\[16\].RFW.BIT\[18\].FF/Q REGF\[16\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[18] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.BIT\[31\].OBUF1 REGF\[17\].RFW.BIT\[31\].FF/Q REGF\[17\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[31] sky130_fd_sc_hd__ebufn_2
Xfill_40_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_40_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[22\].RFW.BIT\[20\].OBUF1 REGF\[22\].RFW.BIT\[20\].FF/Q REGF\[22\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[20] sky130_fd_sc_hd__ebufn_2
Xfill_40_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_49_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_49_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_49_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[7\].RFW.BIT\[10\].OBUF1 REGF\[7\].RFW.BIT\[10\].FF/Q REGF\[7\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[10] sky130_fd_sc_hd__ebufn_2
Xtap_16_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_49_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_49_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[8\].RFW.BIT\[26\].OBUF2 REGF\[8\].RFW.BIT\[26\].FF/Q REGF\[8\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[26] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[21\].OBUF2 REGF\[26\].RFW.BIT\[21\].FF/Q REGF\[26\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[21] sky130_fd_sc_hd__ebufn_2
Xfill_51_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.BIT\[10\].OBUF2 REGF\[31\].RFW.BIT\[10\].FF/Q REGF\[31\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[10] sky130_fd_sc_hd__ebufn_2
Xfill_44_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_37_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_2_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_2_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.BIT\[13\].OBUF1 REGF\[3\].RFW.BIT\[13\].FF/Q REGF\[3\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[13] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.BIT\[29\].OBUF2 REGF\[4\].RFW.BIT\[29\].FF/Q REGF\[4\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[29] sky130_fd_sc_hd__ebufn_2
Xfill_19_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_19_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[22\].RFW.BIT\[24\].OBUF2 REGF\[22\].RFW.BIT\[24\].FF/Q REGF\[22\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[24] sky130_fd_sc_hd__ebufn_2
Xfill_35_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XREGF\[8\].RFW.BIT\[28\].FF REGF\[8\].RFW.CG\[3\]/GCLK DW[28] VGND VGND VPWR VPWR
+ REGF\[8\].RFW.BIT\[28\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[14\].RFW.BIT\[18\].FF REGF\[14\].RFW.CG\[2\]/GCLK DW[18] VGND VGND VPWR VPWR
+ REGF\[14\].RFW.BIT\[18\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[4\].RFW.BIT\[30\].FF REGF\[4\].RFW.CG\[3\]/GCLK DW[30] VGND VGND VPWR VPWR
+ REGF\[4\].RFW.BIT\[30\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[10\].RFW.BIT\[20\].FF REGF\[10\].RFW.CG\[2\]/GCLK DW[20] VGND VGND VPWR VPWR
+ REGF\[10\].RFW.BIT\[20\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_12_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[7\].RFW.BIT\[14\].OBUF2 REGF\[7\].RFW.BIT\[14\].FF/Q REGF\[7\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[14] sky130_fd_sc_hd__ebufn_2
Xfill_51_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_51_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_51_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_51_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.BIT\[22\].OBUF1 REGF\[12\].RFW.BIT\[22\].FF/Q REGF\[12\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[22] sky130_fd_sc_hd__ebufn_2
Xtap_21_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_25_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_25_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[25\].RFW.BIT\[28\].FF REGF\[25\].RFW.CG\[3\]/GCLK DW[28] VGND VGND VPWR VPWR
+ REGF\[25\].RFW.BIT\[28\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[21\].RFW.BIT\[30\].FF REGF\[21\].RFW.CG\[3\]/GCLK DW[30] VGND VGND VPWR VPWR
+ REGF\[21\].RFW.BIT\[30\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_41_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[4\].RFW.BIT\[30\].OBUF2 REGF\[4\].RFW.BIT\[30\].FF/Q REGF\[4\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[30] sky130_fd_sc_hd__ebufn_2
Xgenblk1.RFW0.BIT\[23\].OBUF1 genblk1.RFW0.TIE\[2\]/LO genblk1.RFW0.INV1\[2\]/Y VGND
+ VGND VPWR VPWR DA[23] sky130_fd_sc_hd__ebufn_2
XREGF\[3\].RFW.BIT\[17\].OBUF2 REGF\[3\].RFW.BIT\[17\].FF/Q REGF\[3\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[17] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[23\].OBUF2 REGF\[16\].RFW.BIT\[23\].FF/Q REGF\[16\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[23] sky130_fd_sc_hd__ebufn_2
Xfill_42_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[21\].RFW.BIT\[12\].OBUF2 REGF\[21\].RFW.BIT\[12\].FF/Q REGF\[21\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[12] sky130_fd_sc_hd__ebufn_2
Xfill_35_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_28_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[5\].RFW.BIT\[13\].FF REGF\[5\].RFW.CG\[1\]/GCLK DW[13] VGND VGND VPWR VPWR
+ REGF\[5\].RFW.BIT\[13\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_21_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[11\].RFW.BIT\[10\].OBUF1 REGF\[11\].RFW.BIT\[10\].FF/Q REGF\[11\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[10] sky130_fd_sc_hd__ebufn_2
XDEC0.D0.ABUF\[1\] RA[1] VGND VGND VPWR VPWR DEC0.D0.AND7/B sky130_fd_sc_hd__clkbuf_2
XREGF\[26\].RFW.CG\[1\] CLK REGF\[26\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[26\].RFW.CG\[1\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_46_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_46_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_46_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[12\].RFW.BIT\[26\].OBUF2 REGF\[12\].RFW.BIT\[26\].FF/Q REGF\[12\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[26] sky130_fd_sc_hd__ebufn_2
Xfill_62_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_62_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_62_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[22\].RFW.BIT\[13\].FF REGF\[22\].RFW.CG\[1\]/GCLK DW[13] VGND VGND VPWR VPWR
+ REGF\[22\].RFW.BIT\[13\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_11_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_11_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_11_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[15\].RFW.BIT\[11\].OBUF2 REGF\[15\].RFW.BIT\[11\].FF/Q REGF\[15\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[11] sky130_fd_sc_hd__ebufn_2
XREGF\[7\].RFW.INV2\[2\] DEC1.D0.AND7/X VGND VGND VPWR VPWR REGF\[7\].RFW.INV2\[2\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_21_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgenblk1.RFW0.BIT\[27\].OBUF2 genblk1.RFW0.TIE\[7\]/LO genblk1.RFW0.INV2\[3\]/Y VGND
+ VGND VPWR VPWR DB[27] sky130_fd_sc_hd__ebufn_2
Xfill_14_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[11\].RFW.BIT\[26\].FF REGF\[11\].RFW.CG\[3\]/GCLK DW[26] VGND VGND VPWR VPWR
+ REGF\[11\].RFW.BIT\[26\].FF/Q sky130_fd_sc_hd__dfxtp_1
XDEC2.D2.AND1 DEC2.D2.AND7/C DEC2.D2.AND7/B DEC2.D2.AND7/A DEC2.D2.AND7/D VGND VGND
+ VPWR VPWR DEC2.D2.AND1/X sky130_fd_sc_hd__and4bb_2
XREGF\[17\].RFW.BIT\[20\].FF REGF\[17\].RFW.CG\[2\]/GCLK DW[20] VGND VGND VPWR VPWR
+ REGF\[17\].RFW.BIT\[20\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_8_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[27\].RFW.INV2\[0\] DEC1.D3.AND3/X VGND VGND VPWR VPWR REGF\[27\].RFW.INV2\[0\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_40_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[11\].RFW.BIT\[14\].OBUF2 REGF\[11\].RFW.BIT\[14\].FF/Q REGF\[11\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[14] sky130_fd_sc_hd__ebufn_2
Xfill_16_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[31\].RFW.BIT\[2\].FF REGF\[31\].RFW.CG\[0\]/GCLK DW[2] VGND VGND VPWR VPWR
+ REGF\[31\].RFW.BIT\[2\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[2\].RFW.BIT\[1\].FF REGF\[2\].RFW.CG\[0\]/GCLK DW[1] VGND VGND VPWR VPWR REGF\[2\].RFW.BIT\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[14\].RFW.CG\[1\] CLK REGF\[14\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[14\].RFW.CG\[1\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_32_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_62_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[9\].RFW.BIT\[29\].OBUF1 REGF\[9\].RFW.BIT\[29\].FF/Q REGF\[9\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[29] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.BIT\[30\].FF REGF\[28\].RFW.CG\[3\]/GCLK DW[30] VGND VGND VPWR VPWR
+ REGF\[28\].RFW.BIT\[30\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_48_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.INV1\[3\] DEC0.D0.AND3/X VGND VGND VPWR VPWR REGF\[3\].RFW.INV1\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[27\].RFW.BIT\[24\].OBUF1 REGF\[27\].RFW.BIT\[24\].FF/Q REGF\[27\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[24] sky130_fd_sc_hd__ebufn_2
Xfill_57_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDEC1.D3.AND3 DEC1.D3.AND7/C DEC1.D3.AND7/B DEC1.D3.AND7/A DEC1.D3.AND7/D VGND VGND
+ VPWR VPWR DEC1.D3.AND3/X sky130_fd_sc_hd__and4b_2
Xfill_57_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_57_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_57_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[1\].RFW.BIT\[3\].FF REGF\[1\].RFW.CG\[0\]/GCLK DW[3] VGND VGND VPWR VPWR REGF\[1\].RFW.BIT\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[30\].RFW.BIT\[4\].FF REGF\[30\].RFW.CG\[0\]/GCLK DW[4] VGND VGND VPWR VPWR
+ REGF\[30\].RFW.BIT\[4\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[6\].RFW.BIT\[19\].FF REGF\[6\].RFW.CG\[2\]/GCLK DW[19] VGND VGND VPWR VPWR
+ REGF\[6\].RFW.BIT\[19\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[2\].RFW.BIT\[21\].FF REGF\[2\].RFW.CG\[2\]/GCLK DW[21] VGND VGND VPWR VPWR
+ REGF\[2\].RFW.BIT\[21\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[23\].RFW.INV1\[1\] DEC0.D2.AND7/X VGND VGND VPWR VPWR REGF\[23\].RFW.INV1\[1\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[23\].RFW.BIT\[27\].OBUF1 REGF\[23\].RFW.BIT\[27\].FF/Q REGF\[23\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[27] sky130_fd_sc_hd__ebufn_2
Xfill_12_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[8\].RFW.BIT\[17\].OBUF1 REGF\[8\].RFW.BIT\[17\].FF/Q REGF\[8\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[17] sky130_fd_sc_hd__ebufn_2
XREGF\[23\].RFW.BIT\[19\].FF REGF\[23\].RFW.CG\[2\]/GCLK DW[19] VGND VGND VPWR VPWR
+ REGF\[23\].RFW.BIT\[19\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[9\].RFW.BIT\[30\].OBUF1 REGF\[9\].RFW.BIT\[30\].FF/Q REGF\[9\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[30] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.BIT\[13\].FF REGF\[29\].RFW.CG\[1\]/GCLK DW[13] VGND VGND VPWR VPWR
+ REGF\[29\].RFW.BIT\[13\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[26\].RFW.BIT\[12\].OBUF1 REGF\[26\].RFW.BIT\[12\].FF/Q REGF\[26\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[12] sky130_fd_sc_hd__ebufn_2
Xfill_27_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_27_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_43_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_43_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_43_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XREGF\[27\].RFW.BIT\[28\].OBUF2 REGF\[27\].RFW.BIT\[28\].FF/Q REGF\[27\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[28] sky130_fd_sc_hd__ebufn_2
Xtap_60_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.BIT\[26\].FF REGF\[18\].RFW.CG\[3\]/GCLK DW[26] VGND VGND VPWR VPWR
+ REGF\[18\].RFW.BIT\[26\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_20_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_53_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_46_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[30\].RFW.BIT\[31\].FF REGF\[30\].RFW.CG\[3\]/GCLK DW[31] VGND VGND VPWR VPWR
+ REGF\[30\].RFW.BIT\[31\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_39_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[17\].RFW.BIT\[26\].OBUF1 REGF\[17\].RFW.BIT\[26\].FF/Q REGF\[17\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[26] sky130_fd_sc_hd__ebufn_2
Xfill_17_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_17_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[22\].RFW.BIT\[15\].OBUF1 REGF\[22\].RFW.BIT\[15\].FF/Q REGF\[22\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[15] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.INV1\[2\] DEC0.D2.AND2/X VGND VGND VPWR VPWR REGF\[18\].RFW.INV1\[2\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_33_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_5_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgenblk1.RFW0.TIE\[3\] VGND VGND VPWR VPWR genblk1.RFW0.TIE\[3\]/HI genblk1.RFW0.TIE\[3\]/LO
+ sky130_fd_sc_hd__conb_1
Xfill_5_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_5_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_5_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_10_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_8_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[13\].RFW.BIT\[29\].OBUF1 REGF\[13\].RFW.BIT\[29\].FF/Q REGF\[13\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[29] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[16\].OBUF2 REGF\[26\].RFW.BIT\[16\].FF/Q REGF\[26\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[16] sky130_fd_sc_hd__ebufn_2
XREGF\[3\].RFW.BIT\[27\].FF REGF\[3\].RFW.CG\[3\]/GCLK DW[27] VGND VGND VPWR VPWR
+ REGF\[3\].RFW.BIT\[27\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[9\].RFW.BIT\[21\].FF REGF\[9\].RFW.CG\[2\]/GCLK DW[21] VGND VGND VPWR VPWR
+ REGF\[9\].RFW.BIT\[21\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[15\].RFW.BIT\[11\].FF REGF\[15\].RFW.CG\[1\]/GCLK DW[11] VGND VGND VPWR VPWR
+ REGF\[15\].RFW.BIT\[11\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_32_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[4\].RFW.BIT\[21\].OBUF1 REGF\[4\].RFW.BIT\[21\].FF/Q REGF\[4\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[21] sky130_fd_sc_hd__ebufn_2
XREGF\[31\].RFW.BIT\[14\].FF REGF\[31\].RFW.CG\[1\]/GCLK DW[14] VGND VGND VPWR VPWR
+ REGF\[31\].RFW.BIT\[14\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[16\].RFW.BIT\[14\].OBUF1 REGF\[16\].RFW.BIT\[14\].FF/Q REGF\[16\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[14] sky130_fd_sc_hd__ebufn_2
Xtap_18_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_38_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_38_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_38_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC1.D0.AND6 DEC1.D0.AND7/A DEC1.D0.AND7/B DEC1.D0.AND7/C DEC1.D0.AND7/D VGND VGND
+ VPWR VPWR DEC1.D0.AND6/X sky130_fd_sc_hd__and4b_2
Xfill_54_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_54_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_54_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[27\].FF REGF\[20\].RFW.CG\[3\]/GCLK DW[27] VGND VGND VPWR VPWR
+ REGF\[20\].RFW.BIT\[27\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_51_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[22\].RFW.BIT\[19\].OBUF2 REGF\[22\].RFW.BIT\[19\].FF/Q REGF\[22\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[19] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[21\].FF REGF\[26\].RFW.CG\[2\]/GCLK DW[21] VGND VGND VPWR VPWR
+ REGF\[26\].RFW.BIT\[21\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[8\].RFW.BIT\[22\].OBUF2 REGF\[8\].RFW.BIT\[22\].FF/Q REGF\[8\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[22] sky130_fd_sc_hd__ebufn_2
Xfill_39_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[12\].RFW.BIT\[17\].OBUF1 REGF\[12\].RFW.BIT\[17\].FF/Q REGF\[12\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[17] sky130_fd_sc_hd__ebufn_2
XREGF\[13\].RFW.BIT\[30\].OBUF1 REGF\[13\].RFW.BIT\[30\].FF/Q REGF\[13\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[30] sky130_fd_sc_hd__ebufn_2
XREGF\[12\].RFW.INV2\[3\] DEC1.D1.AND4/X VGND VGND VPWR VPWR REGF\[12\].RFW.INV2\[3\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_58_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_6_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgenblk1.RFW0.BIT\[18\].OBUF1 genblk1.RFW0.TIE\[2\]/LO genblk1.RFW0.INV1\[2\]/Y VGND
+ VGND VPWR VPWR DA[18] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.BIT\[25\].OBUF2 REGF\[4\].RFW.BIT\[25\].FF/Q REGF\[4\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[25] sky130_fd_sc_hd__ebufn_2
Xfill_24_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[5\].RFW.INV1\[0\] DEC0.D0.AND5/X VGND VGND VPWR VPWR REGF\[5\].RFW.INV1\[0\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[16\].RFW.BIT\[18\].OBUF2 REGF\[16\].RFW.BIT\[18\].FF/Q REGF\[16\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[18] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.BIT\[31\].OBUF2 REGF\[17\].RFW.BIT\[31\].FF/Q REGF\[17\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[31] sky130_fd_sc_hd__ebufn_2
Xfill_40_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[22\].RFW.BIT\[20\].OBUF2 REGF\[22\].RFW.BIT\[20\].FF/Q REGF\[22\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[20] sky130_fd_sc_hd__ebufn_2
XDEC1.D3.ABUF\[0\] RB[0] VGND VGND VPWR VPWR DEC1.D3.AND7/A sky130_fd_sc_hd__clkbuf_2
Xtap_30_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_49_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_49_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_49_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[7\].RFW.BIT\[10\].OBUF2 REGF\[7\].RFW.BIT\[10\].FF/Q REGF\[7\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[10] sky130_fd_sc_hd__ebufn_2
Xtap_16_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_49_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_14_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[23\].RFW.CG\[3\] CLK REGF\[23\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[23\].RFW.CG\[3\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[16\].RFW.BIT\[17\].FF REGF\[16\].RFW.CG\[2\]/GCLK DW[17] VGND VGND VPWR VPWR
+ REGF\[16\].RFW.BIT\[17\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_39_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_51_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_44_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_37_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_2_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_2_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_2_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.BIT\[13\].OBUF2 REGF\[3\].RFW.BIT\[13\].FF/Q REGF\[3\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[13] sky130_fd_sc_hd__ebufn_2
XREGF\[22\].RFW.CG\[0\] CLK REGF\[22\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[22\].RFW.CG\[0\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[27\].RFW.BIT\[27\].FF REGF\[27\].RFW.CG\[3\]/GCLK DW[27] VGND VGND VPWR VPWR
+ REGF\[27\].RFW.BIT\[27\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_19_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xtap_12_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_51_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_51_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_51_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XREGF\[1\].RFW.BIT\[18\].FF REGF\[1\].RFW.CG\[2\]/GCLK DW[18] VGND VGND VPWR VPWR
+ REGF\[1\].RFW.BIT\[18\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[12\].RFW.BIT\[22\].OBUF2 REGF\[12\].RFW.BIT\[22\].FF/Q REGF\[12\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[22] sky130_fd_sc_hd__ebufn_2
XREGF\[7\].RFW.BIT\[12\].FF REGF\[7\].RFW.CG\[1\]/GCLK DW[12] VGND VGND VPWR VPWR
+ REGF\[7\].RFW.BIT\[12\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_21_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[11\].RFW.CG\[3\] CLK REGF\[11\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[11\].RFW.CG\[3\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_25_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XREGF\[27\].RFW.BIT\[19\].OBUF1 REGF\[27\].RFW.BIT\[19\].FF/Q REGF\[27\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[19] sky130_fd_sc_hd__ebufn_2
Xfill_41_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_41_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgenblk1.RFW0.BIT\[23\].OBUF2 genblk1.RFW0.TIE\[6\]/LO genblk1.RFW0.INV2\[2\]/Y VGND
+ VGND VPWR VPWR DB[23] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[12\].FF REGF\[24\].RFW.CG\[1\]/GCLK DW[12] VGND VGND VPWR VPWR
+ REGF\[24\].RFW.BIT\[12\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_42_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_28_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XREGF\[10\].RFW.CG\[0\] CLK REGF\[10\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[10\].RFW.CG\[0\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[13\].RFW.BIT\[25\].FF REGF\[13\].RFW.CG\[3\]/GCLK DW[25] VGND VGND VPWR VPWR
+ REGF\[13\].RFW.BIT\[25\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[11\].RFW.BIT\[10\].OBUF2 REGF\[11\].RFW.BIT\[10\].FF/Q REGF\[11\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[10] sky130_fd_sc_hd__ebufn_2
XREGF\[9\].RFW.BIT\[25\].OBUF1 REGF\[9\].RFW.BIT\[25\].FF/Q REGF\[9\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[25] sky130_fd_sc_hd__ebufn_2
Xfill_46_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_0_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_46_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_46_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_62_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_62_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_62_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.INV1\[1\] DEC0.D3.AND7/X VGND VGND VPWR VPWR REGF\[31\].RFW.INV1\[1\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[27\].RFW.BIT\[20\].OBUF1 REGF\[27\].RFW.BIT\[20\].FF/Q REGF\[27\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[20] sky130_fd_sc_hd__ebufn_2
Xfill_11_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_11_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_11_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_11_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XREGF\[14\].RFW.INV2\[0\] DEC1.D1.AND6/X VGND VGND VPWR VPWR REGF\[14\].RFW.INV2\[0\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_21_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_14_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[5\].RFW.BIT\[28\].OBUF1 REGF\[5\].RFW.BIT\[28\].FF/Q REGF\[5\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[28] sky130_fd_sc_hd__ebufn_2
XDEC2.D2.AND2 DEC2.D2.AND7/C DEC2.D2.AND7/A DEC2.D2.AND7/B DEC2.D2.AND7/D VGND VGND
+ VPWR VPWR DEC2.D2.AND2/X sky130_fd_sc_hd__and4bb_2
Xfill_8_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_8_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[23\].RFW.BIT\[23\].OBUF1 REGF\[23\].RFW.BIT\[23\].FF/Q REGF\[23\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[23] sky130_fd_sc_hd__ebufn_2
XREGF\[8\].RFW.BIT\[18\].FF REGF\[8\].RFW.CG\[2\]/GCLK DW[18] VGND VGND VPWR VPWR
+ REGF\[8\].RFW.BIT\[18\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[10\].RFW.BIT\[10\].FF REGF\[10\].RFW.CG\[1\]/GCLK DW[10] VGND VGND VPWR VPWR
+ REGF\[10\].RFW.BIT\[10\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[4\].RFW.BIT\[20\].FF REGF\[4\].RFW.CG\[2\]/GCLK DW[20] VGND VGND VPWR VPWR
+ REGF\[4\].RFW.BIT\[20\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[8\].RFW.BIT\[13\].OBUF1 REGF\[8\].RFW.BIT\[13\].FF/Q REGF\[8\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[13] sky130_fd_sc_hd__ebufn_2
Xfill_40_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_32_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_62_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[9\].RFW.BIT\[29\].OBUF2 REGF\[9\].RFW.BIT\[29\].FF/Q REGF\[9\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[29] sky130_fd_sc_hd__ebufn_2
Xtap_48_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[10\].RFW.INV1\[1\] DEC0.D1.AND2/X VGND VGND VPWR VPWR REGF\[10\].RFW.INV1\[1\]/Y
+ sky130_fd_sc_hd__inv_4
Xtap_18_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[19\].RFW.BIT\[3\].FF REGF\[19\].RFW.CG\[0\]/GCLK DW[3] VGND VGND VPWR VPWR
+ REGF\[19\].RFW.BIT\[3\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[25\].RFW.BIT\[18\].FF REGF\[25\].RFW.CG\[2\]/GCLK DW[18] VGND VGND VPWR VPWR
+ REGF\[25\].RFW.BIT\[18\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_57_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_57_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC1.D3.AND4 DEC1.D3.AND7/A DEC1.D3.AND7/B DEC1.D3.AND7/C DEC1.D3.AND7/D VGND VGND
+ VPWR VPWR DEC1.D3.AND4/X sky130_fd_sc_hd__and4bb_2
XREGF\[27\].RFW.BIT\[24\].OBUF2 REGF\[27\].RFW.BIT\[24\].FF/Q REGF\[27\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[24] sky130_fd_sc_hd__ebufn_2
Xfill_57_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_57_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[21\].RFW.BIT\[20\].FF REGF\[21\].RFW.CG\[2\]/GCLK DW[20] VGND VGND VPWR VPWR
+ REGF\[21\].RFW.BIT\[20\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[26\].RFW.INV1\[2\] DEC0.D3.AND2/X VGND VGND VPWR VPWR REGF\[26\].RFW.INV1\[2\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[4\].RFW.BIT\[16\].OBUF1 REGF\[4\].RFW.BIT\[16\].FF/Q REGF\[4\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[16] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.BIT\[22\].OBUF1 REGF\[17\].RFW.BIT\[22\].FF/Q REGF\[17\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[22] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.BIT\[5\].FF REGF\[18\].RFW.CG\[0\]/GCLK DW[5] VGND VGND VPWR VPWR
+ REGF\[18\].RFW.BIT\[5\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_22_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[22\].RFW.BIT\[11\].OBUF1 REGF\[22\].RFW.BIT\[11\].FF/Q REGF\[22\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[11] sky130_fd_sc_hd__ebufn_2
Xfill_47_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[17\].RFW.BIT\[7\].FF REGF\[17\].RFW.CG\[0\]/GCLK DW[7] VGND VGND VPWR VPWR
+ REGF\[17\].RFW.BIT\[7\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_12_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[23\].RFW.BIT\[27\].OBUF2 REGF\[23\].RFW.BIT\[27\].FF/Q REGF\[23\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[27] sky130_fd_sc_hd__ebufn_2
XREGF\[8\].RFW.BIT\[17\].OBUF2 REGF\[8\].RFW.BIT\[17\].FF/Q REGF\[8\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[17] sky130_fd_sc_hd__ebufn_2
XREGF\[9\].RFW.BIT\[30\].OBUF2 REGF\[9\].RFW.BIT\[30\].FF/Q REGF\[9\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[30] sky130_fd_sc_hd__ebufn_2
XREGF\[13\].RFW.BIT\[25\].OBUF1 REGF\[13\].RFW.BIT\[25\].FF/Q REGF\[13\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[25] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[12\].OBUF2 REGF\[26\].RFW.BIT\[12\].FF/Q REGF\[26\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[12] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[9\].FF REGF\[16\].RFW.CG\[1\]/GCLK DW[9] VGND VGND VPWR VPWR
+ REGF\[16\].RFW.BIT\[9\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_27_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_43_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_43_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[16\].RFW.BIT\[10\].OBUF1 REGF\[16\].RFW.BIT\[10\].FF/Q REGF\[16\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[10] sky130_fd_sc_hd__ebufn_2
Xtap_20_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_60_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_46_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_39_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.CG\[2\] CLK REGF\[31\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[31\].RFW.CG\[2\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[5\].RFW.BIT\[26\].FF REGF\[5\].RFW.CG\[3\]/GCLK DW[26] VGND VGND VPWR VPWR
+ REGF\[5\].RFW.BIT\[26\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[11\].RFW.BIT\[16\].FF REGF\[11\].RFW.CG\[2\]/GCLK DW[16] VGND VGND VPWR VPWR
+ REGF\[11\].RFW.BIT\[16\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[17\].RFW.BIT\[26\].OBUF2 REGF\[17\].RFW.BIT\[26\].FF/Q REGF\[17\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[26] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.BIT\[10\].FF REGF\[17\].RFW.CG\[1\]/GCLK DW[10] VGND VGND VPWR VPWR
+ REGF\[17\].RFW.BIT\[10\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[20\].RFW.INV2\[3\] DEC1.D2.AND4/X VGND VGND VPWR VPWR REGF\[20\].RFW.INV2\[3\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_17_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_17_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[22\].RFW.BIT\[15\].OBUF2 REGF\[22\].RFW.BIT\[15\].FF/Q REGF\[22\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[15] sky130_fd_sc_hd__ebufn_2
Xfill_17_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XREGF\[10\].RFW.BIT\[9\].OBUF1 REGF\[10\].RFW.BIT\[9\].FF/Q REGF\[10\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[9] sky130_fd_sc_hd__ebufn_2
Xfill_33_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[12\].RFW.BIT\[13\].OBUF1 REGF\[12\].RFW.BIT\[13\].FF/Q REGF\[12\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[13] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.BIT\[9\].FF REGF\[29\].RFW.CG\[1\]/GCLK DW[9] VGND VGND VPWR VPWR
+ REGF\[29\].RFW.BIT\[9\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_5_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_5_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_5_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_5_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[22\].RFW.BIT\[26\].FF REGF\[22\].RFW.CG\[3\]/GCLK DW[26] VGND VGND VPWR VPWR
+ REGF\[22\].RFW.BIT\[26\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_5_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[28\].RFW.BIT\[20\].FF REGF\[28\].RFW.CG\[2\]/GCLK DW[20] VGND VGND VPWR VPWR
+ REGF\[28\].RFW.BIT\[20\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_8_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_10_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XREGF\[13\].RFW.BIT\[29\].OBUF2 REGF\[13\].RFW.BIT\[29\].FF/Q REGF\[13\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[29] sky130_fd_sc_hd__ebufn_2
XDEC0.D.AND0 RA[3] RA[4] DEC0.TIE/HI VGND VGND VPWR VPWR DEC0.D.AND0/Y sky130_fd_sc_hd__nor3b_4
Xtap_32_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgenblk1.RFW0.BIT\[14\].OBUF1 genblk1.RFW0.TIE\[1\]/LO genblk1.RFW0.INV1\[1\]/Y VGND
+ VGND VPWR VPWR DA[14] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.BIT\[21\].OBUF2 REGF\[4\].RFW.BIT\[21\].FF/Q REGF\[4\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[21] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[14\].OBUF2 REGF\[16\].RFW.BIT\[14\].FF/Q REGF\[16\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[14] sky130_fd_sc_hd__ebufn_2
Xtap_18_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_38_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDEC1.D0.AND7 DEC1.D0.AND7/A DEC1.D0.AND7/B DEC1.D0.AND7/C DEC1.D0.AND7/D VGND VGND
+ VPWR VPWR DEC1.D0.AND7/X sky130_fd_sc_hd__and4_2
XREGF\[2\].RFW.BIT\[11\].FF REGF\[2\].RFW.CG\[1\]/GCLK DW[11] VGND VGND VPWR VPWR
+ REGF\[2\].RFW.BIT\[11\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[12\].RFW.BIT\[9\].OBUF1 REGF\[12\].RFW.BIT\[9\].FF/Q REGF\[12\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[9] sky130_fd_sc_hd__ebufn_2
Xfill_54_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_54_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_54_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[8\].RFW.CG\[2\] CLK REGF\[8\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[8\].RFW.CG\[2\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_51_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[2\].RFW.BIT\[8\].OBUF1 REGF\[2\].RFW.BIT\[8\].FF/Q REGF\[2\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[8] sky130_fd_sc_hd__ebufn_2
Xtap_44_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.BIT\[17\].OBUF2 REGF\[12\].RFW.BIT\[17\].FF/Q REGF\[12\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[17] sky130_fd_sc_hd__ebufn_2
XREGF\[13\].RFW.BIT\[30\].OBUF2 REGF\[13\].RFW.BIT\[30\].FF/Q REGF\[13\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[30] sky130_fd_sc_hd__ebufn_2
XDEC1.D3.ENBUF DEC1.D.AND3/X VGND VGND VPWR VPWR DEC1.D3.AND7/D sky130_fd_sc_hd__clkbuf_2
XREGF\[14\].RFW.BIT\[9\].OBUF1 REGF\[14\].RFW.BIT\[9\].FF/Q REGF\[14\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[9] sky130_fd_sc_hd__ebufn_2
XREGF\[8\].RFW.INV1\[1\] DEC0.D1.AND0/Y VGND VGND VPWR VPWR REGF\[8\].RFW.INV1\[1\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_58_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[28\].RFW.BIT\[27\].OBUF1 REGF\[28\].RFW.BIT\[27\].FF/Q REGF\[28\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[27] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.BIT\[16\].FF REGF\[18\].RFW.CG\[2\]/GCLK DW[16] VGND VGND VPWR VPWR
+ REGF\[18\].RFW.BIT\[16\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[30\].RFW.BIT\[21\].FF REGF\[30\].RFW.CG\[2\]/GCLK DW[21] VGND VGND VPWR VPWR
+ REGF\[30\].RFW.BIT\[21\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_6_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xgenblk1.RFW0.BIT\[18\].OBUF2 genblk1.RFW0.TIE\[6\]/LO genblk1.RFW0.INV2\[2\]/Y VGND
+ VGND VPWR VPWR DB[18] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.BIT\[8\].OBUF1 REGF\[4\].RFW.BIT\[8\].FF/Q REGF\[4\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[8] sky130_fd_sc_hd__ebufn_2
Xfill_40_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_30_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_23_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_49_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_49_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_49_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xtap_26_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[29\].RFW.BIT\[26\].FF REGF\[29\].RFW.CG\[3\]/GCLK DW[26] VGND VGND VPWR VPWR
+ REGF\[29\].RFW.BIT\[26\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_14_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_14_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[16\].RFW.BIT\[9\].OBUF1 REGF\[16\].RFW.BIT\[9\].FF/Q REGF\[16\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[9] sky130_fd_sc_hd__ebufn_2
Xfill_30_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[27\].RFW.BIT\[15\].OBUF1 REGF\[27\].RFW.BIT\[15\].FF/Q REGF\[27\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[15] sky130_fd_sc_hd__ebufn_2
Xfill_39_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_51_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_44_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.BIT\[17\].FF REGF\[3\].RFW.CG\[2\]/GCLK DW[17] VGND VGND VPWR VPWR
+ REGF\[3\].RFW.BIT\[17\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[6\].RFW.BIT\[8\].OBUF1 REGF\[6\].RFW.BIT\[8\].FF/Q REGF\[6\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[8] sky130_fd_sc_hd__ebufn_2
Xfill_37_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_2_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_2_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_2_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[9\].RFW.BIT\[11\].FF REGF\[9\].RFW.CG\[1\]/GCLK DW[11] VGND VGND VPWR VPWR
+ REGF\[9\].RFW.BIT\[11\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_55_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[14\].RFW.BIT\[0\].FF REGF\[14\].RFW.CG\[0\]/GCLK DW[0] VGND VGND VPWR VPWR
+ REGF\[14\].RFW.BIT\[0\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[2\].RFW.INV2\[2\] DEC1.D0.AND2/X VGND VGND VPWR VPWR REGF\[2\].RFW.INV2\[2\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[18\].RFW.BIT\[29\].OBUF1 REGF\[18\].RFW.BIT\[29\].FF/Q REGF\[18\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[29] sky130_fd_sc_hd__ebufn_2
XREGF\[20\].RFW.BIT\[17\].FF REGF\[20\].RFW.CG\[2\]/GCLK DW[17] VGND VGND VPWR VPWR
+ REGF\[20\].RFW.BIT\[17\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[18\].RFW.BIT\[9\].OBUF1 REGF\[18\].RFW.BIT\[9\].FF/Q REGF\[18\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[9] sky130_fd_sc_hd__ebufn_2
Xfill_35_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[23\].RFW.BIT\[18\].OBUF1 REGF\[23\].RFW.BIT\[18\].FF/Q REGF\[23\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[18] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[31\].OBUF1 REGF\[24\].RFW.BIT\[31\].FF/Q REGF\[24\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[31] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[11\].FF REGF\[26\].RFW.CG\[1\]/GCLK DW[11] VGND VGND VPWR VPWR
+ REGF\[26\].RFW.BIT\[11\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_12_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_51_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[13\].RFW.BIT\[2\].FF REGF\[13\].RFW.CG\[0\]/GCLK DW[2] VGND VGND VPWR VPWR
+ REGF\[13\].RFW.BIT\[2\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_51_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[9\].RFW.BIT\[21\].OBUF1 REGF\[9\].RFW.BIT\[21\].FF/Q REGF\[9\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[21] sky130_fd_sc_hd__ebufn_2
XREGF\[8\].RFW.BIT\[8\].OBUF1 REGF\[8\].RFW.BIT\[8\].FF/Q REGF\[8\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[8] sky130_fd_sc_hd__ebufn_2
XREGF\[22\].RFW.INV2\[0\] DEC1.D2.AND6/X VGND VGND VPWR VPWR REGF\[22\].RFW.INV2\[0\]/Y
+ sky130_fd_sc_hd__inv_4
Xtap_21_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[11\].RFW.BIT\[7\].OBUF1 REGF\[11\].RFW.BIT\[7\].FF/Q REGF\[11\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[7] sky130_fd_sc_hd__ebufn_2
XREGF\[15\].RFW.BIT\[24\].FF REGF\[15\].RFW.CG\[3\]/GCLK DW[24] VGND VGND VPWR VPWR
+ REGF\[15\].RFW.BIT\[24\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[12\].RFW.BIT\[4\].FF REGF\[12\].RFW.CG\[0\]/GCLK DW[4] VGND VGND VPWR VPWR
+ REGF\[12\].RFW.BIT\[4\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_7_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.BIT\[27\].FF REGF\[31\].RFW.CG\[3\]/GCLK DW[27] VGND VGND VPWR VPWR
+ REGF\[31\].RFW.BIT\[27\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_25_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_25_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_25_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[27\].RFW.BIT\[19\].OBUF2 REGF\[27\].RFW.BIT\[19\].FF/Q REGF\[27\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[19] sky130_fd_sc_hd__ebufn_2
Xfill_41_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_41_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[1\].RFW.BIT\[6\].OBUF1 REGF\[1\].RFW.BIT\[6\].FF/Q REGF\[1\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[6] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[0\].FF REGF\[27\].RFW.CG\[0\]/GCLK DW[0] VGND VGND VPWR VPWR
+ REGF\[27\].RFW.BIT\[0\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_41_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[11\].RFW.BIT\[6\].FF REGF\[11\].RFW.CG\[0\]/GCLK DW[6] VGND VGND VPWR VPWR
+ REGF\[11\].RFW.BIT\[6\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[5\].RFW.BIT\[24\].OBUF1 REGF\[5\].RFW.BIT\[24\].FF/Q REGF\[5\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[24] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.BIT\[17\].OBUF1 REGF\[17\].RFW.BIT\[17\].FF/Q REGF\[17\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[17] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.BIT\[30\].OBUF1 REGF\[18\].RFW.BIT\[30\].FF/Q REGF\[18\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[30] sky130_fd_sc_hd__ebufn_2
Xfill_42_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_35_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_28_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[26\].RFW.BIT\[2\].FF REGF\[26\].RFW.CG\[0\]/GCLK DW[2] VGND VGND VPWR VPWR
+ REGF\[26\].RFW.BIT\[2\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[10\].RFW.BIT\[8\].FF REGF\[10\].RFW.CG\[1\]/GCLK DW[8] VGND VGND VPWR VPWR
+ REGF\[10\].RFW.BIT\[8\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[13\].RFW.BIT\[7\].OBUF1 REGF\[13\].RFW.BIT\[7\].FF/Q REGF\[13\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[7] sky130_fd_sc_hd__ebufn_2
XREGF\[25\].RFW.BIT\[4\].FF REGF\[25\].RFW.CG\[0\]/GCLK DW[4] VGND VGND VPWR VPWR
+ REGF\[25\].RFW.BIT\[4\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[9\].RFW.BIT\[25\].OBUF2 REGF\[9\].RFW.BIT\[25\].FF/Q REGF\[9\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[25] sky130_fd_sc_hd__ebufn_2
Xtap_0_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_46_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[1\].RFW.BIT\[27\].OBUF1 REGF\[1\].RFW.BIT\[27\].FF/Q REGF\[1\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[27] sky130_fd_sc_hd__ebufn_2
Xfill_62_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_62_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[3\].RFW.BIT\[6\].OBUF1 REGF\[3\].RFW.BIT\[6\].FF/Q REGF\[3\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[6] sky130_fd_sc_hd__ebufn_2
Xfill_62_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[27\].RFW.BIT\[20\].OBUF2 REGF\[27\].RFW.BIT\[20\].FF/Q REGF\[27\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[20] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.INV2\[1\] DEC1.D2.AND1/X VGND VGND VPWR VPWR REGF\[17\].RFW.INV2\[1\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_11_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_11_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_11_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_11_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_11_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[24\].RFW.BIT\[6\].FF REGF\[24\].RFW.CG\[0\]/GCLK DW[6] VGND VGND VPWR VPWR
+ REGF\[24\].RFW.BIT\[6\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[4\].RFW.BIT\[12\].OBUF1 REGF\[4\].RFW.BIT\[12\].FF/Q REGF\[4\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[12] sky130_fd_sc_hd__ebufn_2
Xfill_36_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_14_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[27\].RFW.BIT\[17\].FF REGF\[27\].RFW.CG\[2\]/GCLK DW[17] VGND VGND VPWR VPWR
+ REGF\[27\].RFW.BIT\[17\].FF/Q sky130_fd_sc_hd__dfxtp_1
XDEC2.D2.AND3 DEC2.D2.AND7/C DEC2.D2.AND7/B DEC2.D2.AND7/A DEC2.D2.AND7/D VGND VGND
+ VPWR VPWR DEC2.D2.AND3/X sky130_fd_sc_hd__and4b_2
XREGF\[23\].RFW.BIT\[8\].FF REGF\[23\].RFW.CG\[1\]/GCLK DW[8] VGND VGND VPWR VPWR
+ REGF\[23\].RFW.BIT\[8\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[5\].RFW.BIT\[28\].OBUF2 REGF\[5\].RFW.BIT\[28\].FF/Q REGF\[5\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[28] sky130_fd_sc_hd__ebufn_2
XREGF\[15\].RFW.BIT\[7\].OBUF1 REGF\[15\].RFW.BIT\[7\].FF/Q REGF\[15\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[7] sky130_fd_sc_hd__ebufn_2
XDEC0.D2.ABUF\[0\] RA[0] VGND VGND VPWR VPWR DEC0.D2.AND7/A sky130_fd_sc_hd__clkbuf_2
Xfill_8_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_8_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_8_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[23\].RFW.BIT\[23\].OBUF2 REGF\[23\].RFW.BIT\[23\].FF/Q REGF\[23\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[23] sky130_fd_sc_hd__ebufn_2
XREGF\[9\].RFW.BIT\[3\].FF REGF\[9\].RFW.CG\[0\]/GCLK DW[3] VGND VGND VPWR VPWR REGF\[9\].RFW.BIT\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[8\].RFW.BIT\[13\].OBUF2 REGF\[8\].RFW.BIT\[13\].FF/Q REGF\[8\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[13] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[6\].OBUF1 REGF\[5\].RFW.BIT\[6\].FF/Q REGF\[5\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[6] sky130_fd_sc_hd__ebufn_2
Xfill_40_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[13\].RFW.INV1\[2\] DEC0.D1.AND5/X VGND VGND VPWR VPWR REGF\[13\].RFW.INV1\[2\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_26_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[13\].RFW.BIT\[21\].OBUF1 REGF\[13\].RFW.BIT\[21\].FF/Q REGF\[13\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[21] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.INV1\[3\] DEC0.D3.AND5/X VGND VGND VPWR VPWR REGF\[29\].RFW.INV1\[3\]/Y
+ sky130_fd_sc_hd__inv_4
Xtap_62_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[8\].RFW.BIT\[5\].FF REGF\[8\].RFW.CG\[0\]/GCLK DW[5] VGND VGND VPWR VPWR REGF\[8\].RFW.BIT\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xtap_48_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_57_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_57_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_57_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC1.D3.AND5 DEC1.D3.AND7/B DEC1.D3.AND7/A DEC1.D3.AND7/C DEC1.D3.AND7/D VGND VGND
+ VPWR VPWR DEC1.D3.AND5/X sky130_fd_sc_hd__and4b_2
XREGF\[17\].RFW.BIT\[7\].OBUF1 REGF\[17\].RFW.BIT\[7\].FF/Q REGF\[17\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[7] sky130_fd_sc_hd__ebufn_2
Xtap_34_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[7\].RFW.BIT\[7\].FF REGF\[7\].RFW.CG\[0\]/GCLK DW[7] VGND VGND VPWR VPWR REGF\[7\].RFW.BIT\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[4\].RFW.BIT\[16\].OBUF2 REGF\[4\].RFW.BIT\[16\].FF/Q REGF\[4\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[16] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.BIT\[22\].OBUF2 REGF\[17\].RFW.BIT\[22\].FF/Q REGF\[17\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[22] sky130_fd_sc_hd__ebufn_2
Xfill_22_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_22_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[7\].RFW.BIT\[6\].OBUF1 REGF\[7\].RFW.BIT\[6\].FF/Q REGF\[7\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[6] sky130_fd_sc_hd__ebufn_2
XREGF\[22\].RFW.BIT\[11\].OBUF2 REGF\[22\].RFW.BIT\[11\].FF/Q REGF\[22\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[11] sky130_fd_sc_hd__ebufn_2
XREGF\[6\].RFW.BIT\[9\].FF REGF\[6\].RFW.CG\[1\]/GCLK DW[9] VGND VGND VPWR VPWR REGF\[6\].RFW.BIT\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[10\].RFW.BIT\[5\].OBUF1 REGF\[10\].RFW.BIT\[5\].FF/Q REGF\[10\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[5] sky130_fd_sc_hd__ebufn_2
Xfill_47_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_47_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[7\].RFW.BIT\[25\].FF REGF\[7\].RFW.CG\[3\]/GCLK DW[25] VGND VGND VPWR VPWR
+ REGF\[7\].RFW.BIT\[25\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_12_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[13\].RFW.BIT\[15\].FF REGF\[13\].RFW.CG\[1\]/GCLK DW[15] VGND VGND VPWR VPWR
+ REGF\[13\].RFW.BIT\[15\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[19\].RFW.BIT\[7\].OBUF1 REGF\[19\].RFW.BIT\[7\].FF/Q REGF\[19\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[7] sky130_fd_sc_hd__ebufn_2
XREGF\[13\].RFW.BIT\[25\].OBUF2 REGF\[13\].RFW.BIT\[25\].FF/Q REGF\[13\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[25] sky130_fd_sc_hd__ebufn_2
Xgenblk1.RFW0.BIT\[10\].OBUF1 genblk1.RFW0.TIE\[1\]/LO genblk1.RFW0.INV1\[1\]/Y VGND
+ VGND VPWR VPWR DA[10] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.CG\[1\] CLK REGF\[4\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[4\].RFW.CG\[1\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[9\].RFW.BIT\[6\].OBUF1 REGF\[9\].RFW.BIT\[6\].FF/Q REGF\[9\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[6] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[25\].FF REGF\[24\].RFW.CG\[3\]/GCLK DW[25] VGND VGND VPWR VPWR
+ REGF\[24\].RFW.BIT\[25\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_43_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[16\].RFW.BIT\[10\].OBUF2 REGF\[16\].RFW.BIT\[10\].FF/Q REGF\[16\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[10] sky130_fd_sc_hd__ebufn_2
Xtap_60_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_20_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.BIT\[5\].OBUF1 REGF\[12\].RFW.BIT\[5\].FF/Q REGF\[12\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[5] sky130_fd_sc_hd__ebufn_2
Xtap_46_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_39_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_17_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_17_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_17_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_17_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[2\].RFW.BIT\[4\].OBUF1 REGF\[2\].RFW.BIT\[4\].FF/Q REGF\[2\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[4] sky130_fd_sc_hd__ebufn_2
Xfill_33_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[4\].RFW.BIT\[10\].FF REGF\[4\].RFW.CG\[1\]/GCLK DW[10] VGND VGND VPWR VPWR
+ REGF\[4\].RFW.BIT\[10\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[10\].RFW.BIT\[9\].OBUF2 REGF\[10\].RFW.BIT\[9\].FF/Q REGF\[10\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[9] sky130_fd_sc_hd__ebufn_2
Xfill_33_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[12\].RFW.BIT\[13\].OBUF2 REGF\[12\].RFW.BIT\[13\].FF/Q REGF\[12\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[13] sky130_fd_sc_hd__ebufn_2
Xfill_5_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_5_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_5_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_5_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[30\].RFW.BIT\[27\].OBUF1 REGF\[30\].RFW.BIT\[27\].FF/Q REGF\[30\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[27] sky130_fd_sc_hd__ebufn_2
Xfill_8_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_10_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[14\].RFW.BIT\[5\].OBUF1 REGF\[14\].RFW.BIT\[5\].FF/Q REGF\[14\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[5] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.CG\[3\] CLK REGF\[19\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[19\].RFW.CG\[3\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[21\].RFW.BIT\[10\].FF REGF\[21\].RFW.CG\[1\]/GCLK DW[10] VGND VGND VPWR VPWR
+ REGF\[21\].RFW.BIT\[10\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[28\].RFW.BIT\[23\].OBUF1 REGF\[28\].RFW.BIT\[23\].FF/Q REGF\[28\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[23] sky130_fd_sc_hd__ebufn_2
XDEC0.D.AND1 RA[4] RA[3] DEC0.TIE/HI VGND VGND VPWR VPWR DEC0.D.AND1/X sky130_fd_sc_hd__and3b_4
Xgenblk1.RFW0.BIT\[14\].OBUF2 genblk1.RFW0.TIE\[5\]/LO genblk1.RFW0.INV2\[1\]/Y VGND
+ VGND VPWR VPWR DB[14] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.BIT\[4\].OBUF1 REGF\[4\].RFW.BIT\[4\].FF/Q REGF\[4\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[4] sky130_fd_sc_hd__ebufn_2
Xtap_18_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_38_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.BIT\[9\].OBUF2 REGF\[12\].RFW.BIT\[9\].FF/Q REGF\[12\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[9] sky130_fd_sc_hd__ebufn_2
Xfill_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_54_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[10\].RFW.BIT\[23\].FF REGF\[10\].RFW.CG\[2\]/GCLK DW[23] VGND VGND VPWR VPWR
+ REGF\[10\].RFW.BIT\[23\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[18\].RFW.CG\[0\] CLK REGF\[18\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[18\].RFW.CG\[0\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_51_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[2\].RFW.BIT\[8\].OBUF2 REGF\[2\].RFW.BIT\[8\].FF/Q REGF\[2\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[8] sky130_fd_sc_hd__ebufn_2
Xtap_44_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_37_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[24\].RFW.BIT\[26\].OBUF1 REGF\[24\].RFW.BIT\[26\].FF/Q REGF\[24\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[26] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[5\].OBUF1 REGF\[16\].RFW.BIT\[5\].FF/Q REGF\[16\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[5] sky130_fd_sc_hd__ebufn_2
Xfill_28_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[9\].RFW.BIT\[16\].OBUF1 REGF\[9\].RFW.BIT\[16\].FF/Q REGF\[9\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[16] sky130_fd_sc_hd__ebufn_2
Xfill_44_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[27\].RFW.BIT\[11\].OBUF1 REGF\[27\].RFW.BIT\[11\].FF/Q REGF\[27\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[11] sky130_fd_sc_hd__ebufn_2
XREGF\[6\].RFW.BIT\[4\].OBUF1 REGF\[6\].RFW.BIT\[4\].FF/Q REGF\[6\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[4] sky130_fd_sc_hd__ebufn_2
XREGF\[14\].RFW.BIT\[9\].OBUF2 REGF\[14\].RFW.BIT\[9\].FF/Q REGF\[14\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[9] sky130_fd_sc_hd__ebufn_2
Xfill_58_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[1\].FF REGF\[20\].RFW.CG\[0\]/GCLK DW[1] VGND VGND VPWR VPWR
+ REGF\[20\].RFW.BIT\[1\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[28\].RFW.BIT\[27\].OBUF2 REGF\[28\].RFW.BIT\[27\].FF/Q REGF\[28\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[27] sky130_fd_sc_hd__ebufn_2
XREGF\[20\].RFW.BIT\[29\].OBUF1 REGF\[20\].RFW.BIT\[29\].FF/Q REGF\[20\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[29] sky130_fd_sc_hd__ebufn_2
Xfill_6_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XREGF\[4\].RFW.BIT\[8\].OBUF2 REGF\[4\].RFW.BIT\[8\].FF/Q REGF\[4\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[8] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[16\].FF REGF\[5\].RFW.CG\[2\]/GCLK DW[16] VGND VGND VPWR VPWR
+ REGF\[5\].RFW.BIT\[16\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[5\].RFW.BIT\[19\].OBUF1 REGF\[5\].RFW.BIT\[19\].FF/Q REGF\[5\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[19] sky130_fd_sc_hd__ebufn_2
XREGF\[30\].RFW.INV2\[0\] DEC1.D3.AND6/X VGND VGND VPWR VPWR REGF\[30\].RFW.INV2\[0\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[18\].RFW.BIT\[25\].OBUF1 REGF\[18\].RFW.BIT\[25\].FF/Q REGF\[18\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[25] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.BIT\[5\].OBUF1 REGF\[18\].RFW.BIT\[5\].FF/Q REGF\[18\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[5] sky130_fd_sc_hd__ebufn_2
Xtap_30_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[23\].RFW.BIT\[14\].OBUF1 REGF\[23\].RFW.BIT\[14\].FF/Q REGF\[23\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[14] sky130_fd_sc_hd__ebufn_2
Xfill_49_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_49_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xtap_16_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[8\].RFW.BIT\[4\].OBUF1 REGF\[8\].RFW.BIT\[4\].FF/Q REGF\[8\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[4] sky130_fd_sc_hd__ebufn_2
Xtap_42_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_14_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_14_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_14_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[22\].RFW.BIT\[16\].FF REGF\[22\].RFW.CG\[2\]/GCLK DW[16] VGND VGND VPWR VPWR
+ REGF\[22\].RFW.BIT\[16\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[16\].RFW.BIT\[9\].OBUF2 REGF\[16\].RFW.BIT\[9\].FF/Q REGF\[16\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[9] sky130_fd_sc_hd__ebufn_2
XREGF\[11\].RFW.BIT\[3\].OBUF1 REGF\[11\].RFW.BIT\[3\].FF/Q REGF\[11\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[3] sky130_fd_sc_hd__ebufn_2
Xfill_30_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_30_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[28\].RFW.BIT\[10\].FF REGF\[28\].RFW.CG\[1\]/GCLK DW[10] VGND VGND VPWR VPWR
+ REGF\[28\].RFW.BIT\[10\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[4\].RFW.BIT\[0\].FF REGF\[4\].RFW.CG\[0\]/GCLK DW[0] VGND VGND VPWR VPWR REGF\[4\].RFW.BIT\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[14\].RFW.BIT\[28\].OBUF1 REGF\[14\].RFW.BIT\[28\].FF/Q REGF\[14\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[28] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[15\].OBUF2 REGF\[27\].RFW.BIT\[15\].FF/Q REGF\[27\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[15] sky130_fd_sc_hd__ebufn_2
Xfill_39_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_44_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.BIT\[8\].OBUF2 REGF\[6\].RFW.BIT\[8\].FF/Q REGF\[6\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[8] sky130_fd_sc_hd__ebufn_2
XREGF\[1\].RFW.BIT\[2\].OBUF1 REGF\[1\].RFW.BIT\[2\].FF/Q REGF\[1\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[2] sky130_fd_sc_hd__ebufn_2
Xfill_37_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_2_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_2_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[20\].RFW.BIT\[30\].OBUF1 REGF\[20\].RFW.BIT\[30\].FF/Q REGF\[20\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[30] sky130_fd_sc_hd__ebufn_2
Xfill_55_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_55_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[11\].RFW.BIT\[29\].FF REGF\[11\].RFW.CG\[3\]/GCLK DW[29] VGND VGND VPWR VPWR
+ REGF\[11\].RFW.BIT\[29\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_2_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[5\].RFW.BIT\[20\].OBUF1 REGF\[5\].RFW.BIT\[20\].FF/Q REGF\[5\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[20] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.INV2\[3\] DEC1.D0.AND5/X VGND VGND VPWR VPWR REGF\[5\].RFW.INV2\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[17\].RFW.BIT\[23\].FF REGF\[17\].RFW.CG\[2\]/GCLK DW[23] VGND VGND VPWR VPWR
+ REGF\[17\].RFW.BIT\[23\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[17\].RFW.BIT\[13\].OBUF1 REGF\[17\].RFW.BIT\[13\].FF/Q REGF\[17\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[13] sky130_fd_sc_hd__ebufn_2
XREGF\[3\].RFW.BIT\[2\].FF REGF\[3\].RFW.CG\[0\]/GCLK DW[2] VGND VGND VPWR VPWR REGF\[3\].RFW.BIT\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xfill_56_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.BIT\[29\].OBUF2 REGF\[18\].RFW.BIT\[29\].FF/Q REGF\[18\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[29] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.BIT\[9\].OBUF2 REGF\[18\].RFW.BIT\[9\].FF/Q REGF\[18\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[9] sky130_fd_sc_hd__ebufn_2
XREGF\[25\].RFW.INV2\[1\] DEC1.D3.AND1/X VGND VGND VPWR VPWR REGF\[25\].RFW.INV2\[1\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[31\].RFW.BIT\[5\].FF REGF\[31\].RFW.CG\[0\]/GCLK DW[5] VGND VGND VPWR VPWR
+ REGF\[31\].RFW.BIT\[5\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[13\].RFW.BIT\[3\].OBUF1 REGF\[13\].RFW.BIT\[3\].FF/Q REGF\[13\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[3] sky130_fd_sc_hd__ebufn_2
XREGF\[2\].RFW.BIT\[4\].FF REGF\[2\].RFW.CG\[0\]/GCLK DW[4] VGND VGND VPWR VPWR REGF\[2\].RFW.BIT\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[23\].RFW.BIT\[18\].OBUF2 REGF\[23\].RFW.BIT\[18\].FF/Q REGF\[23\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[18] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[31\].OBUF2 REGF\[24\].RFW.BIT\[31\].FF/Q REGF\[24\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[31] sky130_fd_sc_hd__ebufn_2
Xfill_51_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[9\].RFW.BIT\[21\].OBUF2 REGF\[9\].RFW.BIT\[21\].FF/Q REGF\[9\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[21] sky130_fd_sc_hd__ebufn_2
XREGF\[8\].RFW.BIT\[8\].OBUF2 REGF\[8\].RFW.BIT\[8\].FF/Q REGF\[8\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[8] sky130_fd_sc_hd__ebufn_2
XREGF\[1\].RFW.BIT\[23\].OBUF1 REGF\[1\].RFW.BIT\[23\].FF/Q REGF\[1\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[23] sky130_fd_sc_hd__ebufn_2
XREGF\[3\].RFW.BIT\[2\].OBUF1 REGF\[3\].RFW.BIT\[2\].FF/Q REGF\[3\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[2] sky130_fd_sc_hd__ebufn_2
XREGF\[13\].RFW.BIT\[16\].OBUF1 REGF\[13\].RFW.BIT\[16\].FF/Q REGF\[13\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[16] sky130_fd_sc_hd__ebufn_2
Xtap_21_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[1\].RFW.BIT\[6\].FF REGF\[1\].RFW.CG\[0\]/GCLK DW[6] VGND VGND VPWR VPWR REGF\[1\].RFW.BIT\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xtap_14_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[30\].RFW.BIT\[7\].FF REGF\[30\].RFW.CG\[0\]/GCLK DW[7] VGND VGND VPWR VPWR
+ REGF\[30\].RFW.BIT\[7\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[11\].RFW.BIT\[7\].OBUF2 REGF\[11\].RFW.BIT\[7\].FF/Q REGF\[11\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[7] sky130_fd_sc_hd__ebufn_2
Xtap_7_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC1.D2.ENBUF DEC1.D.AND2/X VGND VGND VPWR VPWR DEC1.D2.AND7/D sky130_fd_sc_hd__clkbuf_2
Xfill_25_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_25_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_25_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_25_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XREGF\[2\].RFW.BIT\[24\].FF REGF\[2\].RFW.CG\[3\]/GCLK DW[24] VGND VGND VPWR VPWR
+ REGF\[2\].RFW.BIT\[24\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_41_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_41_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[1\].RFW.BIT\[6\].OBUF2 REGF\[1\].RFW.BIT\[6\].FF/Q REGF\[1\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[6] sky130_fd_sc_hd__ebufn_2
Xfill_41_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_41_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[30\].RFW.BIT\[11\].FF REGF\[30\].RFW.CG\[1\]/GCLK DW[11] VGND VGND VPWR VPWR
+ REGF\[30\].RFW.BIT\[11\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[5\].RFW.BIT\[24\].OBUF2 REGF\[5\].RFW.BIT\[24\].FF/Q REGF\[5\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[24] sky130_fd_sc_hd__ebufn_2
XREGF\[15\].RFW.BIT\[3\].OBUF1 REGF\[15\].RFW.BIT\[3\].FF/Q REGF\[15\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[3] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.INV1\[2\] DEC0.D2.AND5/X VGND VGND VPWR VPWR REGF\[21\].RFW.INV1\[2\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[17\].RFW.BIT\[17\].OBUF2 REGF\[17\].RFW.BIT\[17\].FF/Q REGF\[17\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[17] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.BIT\[30\].OBUF2 REGF\[18\].RFW.BIT\[30\].FF/Q REGF\[18\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[30] sky130_fd_sc_hd__ebufn_2
Xfill_42_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_35_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_28_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[5\].RFW.BIT\[2\].OBUF1 REGF\[5\].RFW.BIT\[2\].FF/Q REGF\[5\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[2] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.BIT\[16\].FF REGF\[29\].RFW.CG\[2\]/GCLK DW[16] VGND VGND VPWR VPWR
+ REGF\[29\].RFW.BIT\[16\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[13\].RFW.BIT\[7\].OBUF2 REGF\[13\].RFW.BIT\[7\].FF/Q REGF\[13\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[7] sky130_fd_sc_hd__ebufn_2
Xtap_0_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_46_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[1\].RFW.BIT\[27\].OBUF2 REGF\[1\].RFW.BIT\[27\].FF/Q REGF\[1\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[27] sky130_fd_sc_hd__ebufn_2
Xfill_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_62_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.BIT\[6\].OBUF2 REGF\[3\].RFW.BIT\[6\].FF/Q REGF\[3\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[6] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.BIT\[29\].FF REGF\[18\].RFW.CG\[3\]/GCLK DW[29] VGND VGND VPWR VPWR
+ REGF\[18\].RFW.BIT\[29\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[14\].RFW.BIT\[31\].FF REGF\[14\].RFW.CG\[3\]/GCLK DW[31] VGND VGND VPWR VPWR
+ REGF\[14\].RFW.BIT\[31\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[17\].RFW.BIT\[3\].OBUF1 REGF\[17\].RFW.BIT\[3\].FF/Q REGF\[17\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[3] sky130_fd_sc_hd__ebufn_2
Xfill_11_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_11_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_11_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_11_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgenblk1.RFW0.BIT\[7\].OBUF1 genblk1.RFW0.TIE\[0\]/LO genblk1.RFW0.INV1\[0\]/Y VGND
+ VGND VPWR VPWR DA[7] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.BIT\[12\].OBUF2 REGF\[4\].RFW.BIT\[12\].FF/Q REGF\[4\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[12] sky130_fd_sc_hd__ebufn_2
XREGF\[1\].RFW.CG\[3\] CLK REGF\[1\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[1\].RFW.CG\[3\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[7\].RFW.BIT\[2\].OBUF1 REGF\[7\].RFW.BIT\[2\].FF/Q REGF\[7\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[2] sky130_fd_sc_hd__ebufn_2
Xfill_36_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_36_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDEC2.D2.AND4 DEC2.D2.AND7/A DEC2.D2.AND7/B DEC2.D2.AND7/C DEC2.D2.AND7/D VGND VGND
+ VPWR VPWR DEC2.D2.AND4/X sky130_fd_sc_hd__and4bb_2
Xfill_52_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[15\].RFW.BIT\[7\].OBUF2 REGF\[15\].RFW.BIT\[7\].FF/Q REGF\[15\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[7] sky130_fd_sc_hd__ebufn_2
XREGF\[10\].RFW.BIT\[1\].OBUF1 REGF\[10\].RFW.BIT\[1\].FF/Q REGF\[10\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[1] sky130_fd_sc_hd__ebufn_2
Xfill_8_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_8_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[27\].RFW.CG\[2\] CLK REGF\[27\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[27\].RFW.CG\[2\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_8_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[16\].RFW.INV1\[3\] DEC0.D2.AND0/Y VGND VGND VPWR VPWR REGF\[16\].RFW.INV1\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[5\].RFW.BIT\[6\].OBUF2 REGF\[5\].RFW.BIT\[6\].FF/Q REGF\[5\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[6] sky130_fd_sc_hd__ebufn_2
Xfill_40_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_26_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_19_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[19\].RFW.BIT\[3\].OBUF1 REGF\[19\].RFW.BIT\[3\].FF/Q REGF\[19\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[3] sky130_fd_sc_hd__ebufn_2
XREGF\[13\].RFW.BIT\[21\].OBUF2 REGF\[13\].RFW.BIT\[21\].FF/Q REGF\[13\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[21] sky130_fd_sc_hd__ebufn_2
XREGF\[9\].RFW.BIT\[24\].FF REGF\[9\].RFW.CG\[3\]/GCLK DW[24] VGND VGND VPWR VPWR
+ REGF\[9\].RFW.BIT\[24\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[15\].RFW.BIT\[14\].FF REGF\[15\].RFW.CG\[1\]/GCLK DW[14] VGND VGND VPWR VPWR
+ REGF\[15\].RFW.BIT\[14\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_48_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.BIT\[17\].FF REGF\[31\].RFW.CG\[2\]/GCLK DW[17] VGND VGND VPWR VPWR
+ REGF\[31\].RFW.BIT\[17\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[9\].RFW.BIT\[2\].OBUF1 REGF\[9\].RFW.BIT\[2\].FF/Q REGF\[9\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[2] sky130_fd_sc_hd__ebufn_2
Xfill_57_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_18_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_57_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDEC1.D3.AND6 DEC1.D3.AND7/A DEC1.D3.AND7/B DEC1.D3.AND7/C DEC1.D3.AND7/D VGND VGND
+ VPWR VPWR DEC1.D3.AND6/X sky130_fd_sc_hd__and4b_2
XREGF\[28\].RFW.BIT\[18\].OBUF1 REGF\[28\].RFW.BIT\[18\].FF/Q REGF\[28\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[18] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.BIT\[31\].OBUF1 REGF\[29\].RFW.BIT\[31\].FF/Q REGF\[29\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[31] sky130_fd_sc_hd__ebufn_2
XREGF\[12\].RFW.BIT\[1\].OBUF1 REGF\[12\].RFW.BIT\[1\].FF/Q REGF\[12\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[1] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.BIT\[7\].OBUF2 REGF\[17\].RFW.BIT\[7\].FF/Q REGF\[17\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[7] sky130_fd_sc_hd__ebufn_2
Xtap_34_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_50_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_22_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_22_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_22_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[7\].RFW.BIT\[6\].OBUF2 REGF\[7\].RFW.BIT\[6\].FF/Q REGF\[7\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[6] sky130_fd_sc_hd__ebufn_2
XREGF\[2\].RFW.BIT\[0\].OBUF1 REGF\[2\].RFW.BIT\[0\].FF/Q REGF\[2\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[0] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[24\].FF REGF\[26\].RFW.CG\[3\]/GCLK DW[24] VGND VGND VPWR VPWR
+ REGF\[26\].RFW.BIT\[24\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[10\].RFW.BIT\[5\].OBUF2 REGF\[10\].RFW.BIT\[5\].FF/Q REGF\[10\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[5] sky130_fd_sc_hd__ebufn_2
XREGF\[7\].RFW.INV2\[0\] DEC1.D0.AND7/X VGND VGND VPWR VPWR REGF\[7\].RFW.INV2\[0\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_47_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_47_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_47_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_12_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[15\].RFW.CG\[2\] CLK REGF\[15\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[15\].RFW.CG\[2\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[30\].RFW.BIT\[23\].OBUF1 REGF\[30\].RFW.BIT\[23\].FF/Q REGF\[30\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[23] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.BIT\[7\].OBUF2 REGF\[19\].RFW.BIT\[7\].FF/Q REGF\[19\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[7] sky130_fd_sc_hd__ebufn_2
XREGF\[14\].RFW.BIT\[1\].OBUF1 REGF\[14\].RFW.BIT\[1\].FF/Q REGF\[14\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[1] sky130_fd_sc_hd__ebufn_2
Xgenblk1.RFW0.BIT\[10\].OBUF2 genblk1.RFW0.TIE\[5\]/LO genblk1.RFW0.INV2\[1\]/Y VGND
+ VGND VPWR VPWR DB[10] sky130_fd_sc_hd__ebufn_2
XREGF\[9\].RFW.BIT\[6\].OBUF2 REGF\[9\].RFW.BIT\[6\].FF/Q REGF\[9\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[6] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.BIT\[0\].OBUF1 REGF\[4\].RFW.BIT\[0\].FF/Q REGF\[4\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[0] sky130_fd_sc_hd__ebufn_2
Xtap_60_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.BIT\[5\].OBUF2 REGF\[12\].RFW.BIT\[5\].FF/Q REGF\[12\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[5] sky130_fd_sc_hd__ebufn_2
Xtap_46_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.INV1\[1\] DEC0.D0.AND3/X VGND VGND VPWR VPWR REGF\[3\].RFW.INV1\[1\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[6\].RFW.BIT\[27\].OBUF1 REGF\[6\].RFW.BIT\[27\].FF/Q REGF\[6\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[27] sky130_fd_sc_hd__ebufn_2
Xfill_17_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_17_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_17_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_17_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[2\].RFW.BIT\[4\].OBUF2 REGF\[2\].RFW.BIT\[4\].FF/Q REGF\[2\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[4] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[22\].OBUF1 REGF\[24\].RFW.BIT\[22\].FF/Q REGF\[24\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[22] sky130_fd_sc_hd__ebufn_2
Xfill_33_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[16\].RFW.BIT\[1\].OBUF1 REGF\[16\].RFW.BIT\[1\].FF/Q REGF\[16\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[1] sky130_fd_sc_hd__ebufn_2
Xfill_33_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[9\].RFW.BIT\[12\].OBUF1 REGF\[9\].RFW.BIT\[12\].FF/Q REGF\[9\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[12] sky130_fd_sc_hd__ebufn_2
XREGF\[12\].RFW.BIT\[22\].FF REGF\[12\].RFW.CG\[2\]/GCLK DW[22] VGND VGND VPWR VPWR
+ REGF\[12\].RFW.BIT\[22\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_5_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_5_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_5_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_5_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_5_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[6\].RFW.BIT\[0\].OBUF1 REGF\[6\].RFW.BIT\[0\].FF/Q REGF\[6\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[0] sky130_fd_sc_hd__ebufn_2
XREGF\[30\].RFW.BIT\[27\].OBUF2 REGF\[30\].RFW.BIT\[27\].FF/Q REGF\[30\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[27] sky130_fd_sc_hd__ebufn_2
Xfill_8_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_10_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[14\].RFW.BIT\[5\].OBUF2 REGF\[14\].RFW.BIT\[5\].FF/Q REGF\[14\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[5] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.BIT\[23\].OBUF2 REGF\[28\].RFW.BIT\[23\].FF/Q REGF\[28\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[23] sky130_fd_sc_hd__ebufn_2
XREGF\[20\].RFW.BIT\[25\].OBUF1 REGF\[20\].RFW.BIT\[25\].FF/Q REGF\[20\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[25] sky130_fd_sc_hd__ebufn_2
XDEC0.D.AND2 RA[3] RA[4] DEC0.TIE/HI VGND VGND VPWR VPWR DEC0.D.AND2/X sky130_fd_sc_hd__and3b_4
XREGF\[5\].RFW.BIT\[15\].OBUF1 REGF\[5\].RFW.BIT\[15\].FF/Q REGF\[5\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[15] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.BIT\[4\].OBUF2 REGF\[4\].RFW.BIT\[4\].FF/Q REGF\[4\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[4] sky130_fd_sc_hd__ebufn_2
Xtap_18_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.BIT\[21\].OBUF1 REGF\[18\].RFW.BIT\[21\].FF/Q REGF\[18\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[21] sky130_fd_sc_hd__ebufn_2
Xfill_54_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.BIT\[1\].OBUF1 REGF\[18\].RFW.BIT\[1\].FF/Q REGF\[18\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[1] sky130_fd_sc_hd__ebufn_2
XREGF\[23\].RFW.BIT\[10\].OBUF1 REGF\[23\].RFW.BIT\[10\].FF/Q REGF\[23\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[10] sky130_fd_sc_hd__ebufn_2
Xtap_51_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_44_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[8\].RFW.BIT\[0\].OBUF1 REGF\[8\].RFW.BIT\[0\].FF/Q REGF\[8\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[0] sky130_fd_sc_hd__ebufn_2
XREGF\[7\].RFW.BIT\[15\].FF REGF\[7\].RFW.CG\[1\]/GCLK DW[15] VGND VGND VPWR VPWR
+ REGF\[7\].RFW.BIT\[15\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_37_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[24\].RFW.BIT\[26\].OBUF2 REGF\[24\].RFW.BIT\[26\].FF/Q REGF\[24\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[26] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[5\].OBUF2 REGF\[16\].RFW.BIT\[5\].FF/Q REGF\[16\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[5] sky130_fd_sc_hd__ebufn_2
Xfill_28_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_28_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[9\].RFW.BIT\[16\].OBUF2 REGF\[9\].RFW.BIT\[16\].FF/Q REGF\[9\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[16] sky130_fd_sc_hd__ebufn_2
XREGF\[1\].RFW.BIT\[18\].OBUF1 REGF\[1\].RFW.BIT\[18\].FF/Q REGF\[1\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[18] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.INV1\[0\] DEC0.D2.AND2/X VGND VGND VPWR VPWR REGF\[18\].RFW.INV1\[0\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[2\].RFW.BIT\[31\].OBUF1 REGF\[2\].RFW.BIT\[31\].FF/Q REGF\[2\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[31] sky130_fd_sc_hd__ebufn_2
Xfill_44_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_44_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[14\].RFW.BIT\[24\].OBUF1 REGF\[14\].RFW.BIT\[24\].FF/Q REGF\[14\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[24] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[11\].OBUF2 REGF\[27\].RFW.BIT\[11\].FF/Q REGF\[27\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[11] sky130_fd_sc_hd__ebufn_2
Xfill_60_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[6\].RFW.BIT\[4\].OBUF2 REGF\[6\].RFW.BIT\[4\].FF/Q REGF\[6\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[4] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[15\].FF REGF\[24\].RFW.CG\[1\]/GCLK DW[15] VGND VGND VPWR VPWR
+ REGF\[24\].RFW.BIT\[15\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xgenblk1.RFW0.TIE\[1\] VGND VGND VPWR VPWR genblk1.RFW0.TIE\[1\]/HI genblk1.RFW0.TIE\[1\]/LO
+ sky130_fd_sc_hd__conb_1
Xfill_58_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[29\].OBUF2 REGF\[20\].RFW.BIT\[29\].FF/Q REGF\[20\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[29] sky130_fd_sc_hd__ebufn_2
Xfill_6_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[5\].RFW.BIT\[19\].OBUF2 REGF\[5\].RFW.BIT\[19\].FF/Q REGF\[5\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[19] sky130_fd_sc_hd__ebufn_2
XREGF\[13\].RFW.BIT\[28\].FF REGF\[13\].RFW.CG\[3\]/GCLK DW[28] VGND VGND VPWR VPWR
+ REGF\[13\].RFW.BIT\[28\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[18\].RFW.BIT\[25\].OBUF2 REGF\[18\].RFW.BIT\[25\].FF/Q REGF\[18\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[25] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.BIT\[5\].OBUF2 REGF\[18\].RFW.BIT\[5\].FF/Q REGF\[18\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[5] sky130_fd_sc_hd__ebufn_2
XREGF\[10\].RFW.BIT\[27\].OBUF1 REGF\[10\].RFW.BIT\[27\].FF/Q REGF\[10\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[27] sky130_fd_sc_hd__ebufn_2
Xtap_30_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[23\].RFW.BIT\[14\].OBUF2 REGF\[23\].RFW.BIT\[14\].FF/Q REGF\[23\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[14] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.BIT\[22\].FF REGF\[19\].RFW.CG\[2\]/GCLK DW[22] VGND VGND VPWR VPWR
+ REGF\[19\].RFW.BIT\[22\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_49_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_9_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[8\].OBUF1 REGF\[20\].RFW.BIT\[8\].FF/Q REGF\[20\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[8] sky130_fd_sc_hd__ebufn_2
XREGF\[8\].RFW.BIT\[4\].OBUF2 REGF\[8\].RFW.BIT\[4\].FF/Q REGF\[8\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[4] sky130_fd_sc_hd__ebufn_2
Xtap_42_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[13\].RFW.BIT\[12\].OBUF1 REGF\[13\].RFW.BIT\[12\].FF/Q REGF\[13\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[12] sky130_fd_sc_hd__ebufn_2
Xfill_14_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_14_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_14_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[11\].RFW.BIT\[3\].OBUF2 REGF\[11\].RFW.BIT\[3\].FF/Q REGF\[11\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[3] sky130_fd_sc_hd__ebufn_2
XREGF\[9\].RFW.CGAND DEC2.D1.AND1/X WE VGND VGND VPWR VPWR REGF\[9\].RFW.CGAND/X sky130_fd_sc_hd__and2_1
Xfill_30_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_30_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_30_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC0.D0.AND0 DEC0.D0.AND7/A DEC0.D0.AND7/B DEC0.D0.AND7/C DEC0.D0.AND7/D VGND VGND
+ VPWR VPWR DEC0.D0.AND0/Y sky130_fd_sc_hd__nor4b_2
XREGF\[14\].RFW.BIT\[28\].OBUF2 REGF\[14\].RFW.BIT\[28\].FF/Q REGF\[14\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[28] sky130_fd_sc_hd__ebufn_2
Xfill_39_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_39_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_37_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_2_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[1\].RFW.BIT\[2\].OBUF2 REGF\[1\].RFW.BIT\[2\].FF/Q REGF\[1\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[2] sky130_fd_sc_hd__ebufn_2
Xfill_2_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[30\].OBUF2 REGF\[20\].RFW.BIT\[30\].FF/Q REGF\[20\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[30] sky130_fd_sc_hd__ebufn_2
Xfill_55_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_55_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_55_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_2_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[5\].RFW.BIT\[20\].OBUF2 REGF\[5\].RFW.BIT\[20\].FF/Q REGF\[5\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[20] sky130_fd_sc_hd__ebufn_2
XREGF\[12\].RFW.INV2\[1\] DEC1.D1.AND4/X VGND VGND VPWR VPWR REGF\[12\].RFW.INV2\[1\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[17\].RFW.BIT\[13\].OBUF2 REGF\[17\].RFW.BIT\[13\].FF/Q REGF\[17\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[13] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.INV2\[2\] DEC1.D3.AND4/X VGND VGND VPWR VPWR REGF\[28\].RFW.INV2\[2\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[22\].RFW.BIT\[8\].OBUF1 REGF\[22\].RFW.BIT\[8\].FF/Q REGF\[22\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[8] sky130_fd_sc_hd__ebufn_2
XREGF\[10\].RFW.BIT\[13\].FF REGF\[10\].RFW.CG\[1\]/GCLK DW[13] VGND VGND VPWR VPWR
+ REGF\[10\].RFW.BIT\[13\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[4\].RFW.BIT\[23\].FF REGF\[4\].RFW.CG\[2\]/GCLK DW[23] VGND VGND VPWR VPWR
+ REGF\[4\].RFW.BIT\[23\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_56_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_49_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[13\].RFW.BIT\[3\].OBUF2 REGF\[13\].RFW.BIT\[3\].FF/Q REGF\[13\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[3] sky130_fd_sc_hd__ebufn_2
Xfill_4_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[1\].RFW.BIT\[23\].OBUF2 REGF\[1\].RFW.BIT\[23\].FF/Q REGF\[1\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[23] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.BIT\[6\].FF REGF\[19\].RFW.CG\[0\]/GCLK DW[6] VGND VGND VPWR VPWR
+ REGF\[19\].RFW.BIT\[6\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[3\].RFW.BIT\[2\].OBUF2 REGF\[3\].RFW.BIT\[2\].FF/Q REGF\[3\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[2] sky130_fd_sc_hd__ebufn_2
Xtap_21_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[13\].RFW.BIT\[16\].OBUF2 REGF\[13\].RFW.BIT\[16\].FF/Q REGF\[13\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[16] sky130_fd_sc_hd__ebufn_2
Xtap_14_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[21\].RFW.BIT\[23\].FF REGF\[21\].RFW.CG\[2\]/GCLK DW[23] VGND VGND VPWR VPWR
+ REGF\[21\].RFW.BIT\[23\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_7_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgenblk1.RFW0.BIT\[3\].OBUF1 genblk1.RFW0.TIE\[0\]/LO genblk1.RFW0.INV1\[0\]/Y VGND
+ VGND VPWR VPWR DA[3] sky130_fd_sc_hd__ebufn_2
Xfill_25_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_25_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_25_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_25_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_25_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[24\].RFW.INV1\[3\] DEC0.D3.AND0/Y VGND VGND VPWR VPWR REGF\[24\].RFW.INV1\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[24\].RFW.BIT\[8\].OBUF1 REGF\[24\].RFW.BIT\[8\].FF/Q REGF\[24\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[8] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.BIT\[8\].FF REGF\[18\].RFW.CG\[1\]/GCLK DW[8] VGND VGND VPWR VPWR
+ REGF\[18\].RFW.BIT\[8\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[23\].RFW.CG\[1\] CLK REGF\[23\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[23\].RFW.CG\[1\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_41_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_41_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_41_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[29\].RFW.BIT\[26\].OBUF1 REGF\[29\].RFW.BIT\[26\].FF/Q REGF\[29\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[26] sky130_fd_sc_hd__ebufn_2
Xfill_41_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_41_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[15\].RFW.BIT\[3\].OBUF2 REGF\[15\].RFW.BIT\[3\].FF/Q REGF\[15\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[3] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[30\].FF REGF\[16\].RFW.CG\[3\]/GCLK DW[30] VGND VGND VPWR VPWR
+ REGF\[16\].RFW.BIT\[30\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_42_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_35_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_28_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[19\].RFW.CGAND DEC2.D2.AND3/X WE VGND VGND VPWR VPWR REGF\[19\].RFW.CGAND/X
+ sky130_fd_sc_hd__and2_1
XREGF\[5\].RFW.BIT\[2\].OBUF2 REGF\[5\].RFW.BIT\[2\].FF/Q REGF\[5\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[2] sky130_fd_sc_hd__ebufn_2
XREGF\[25\].RFW.BIT\[29\].OBUF1 REGF\[25\].RFW.BIT\[29\].FF/Q REGF\[25\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[29] sky130_fd_sc_hd__ebufn_2
Xtap_0_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[26\].RFW.BIT\[8\].OBUF1 REGF\[26\].RFW.BIT\[8\].FF/Q REGF\[26\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[8] sky130_fd_sc_hd__ebufn_2
XREGF\[30\].RFW.BIT\[18\].OBUF1 REGF\[30\].RFW.BIT\[18\].FF/Q REGF\[30\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[18] sky130_fd_sc_hd__ebufn_2
XREGF\[31\].RFW.BIT\[31\].OBUF1 REGF\[31\].RFW.BIT\[31\].FF/Q REGF\[31\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[31] sky130_fd_sc_hd__ebufn_2
Xfill_62_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[28\].RFW.BIT\[14\].OBUF1 REGF\[28\].RFW.BIT\[14\].FF/Q REGF\[28\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[14] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.BIT\[3\].OBUF2 REGF\[17\].RFW.BIT\[3\].FF/Q REGF\[17\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[3] sky130_fd_sc_hd__ebufn_2
Xfill_11_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_11_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_11_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_11_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_11_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgenblk1.RFW0.BIT\[7\].OBUF2 genblk1.RFW0.TIE\[4\]/LO genblk1.RFW0.INV2\[0\]/Y VGND
+ VGND VPWR VPWR DB[7] sky130_fd_sc_hd__ebufn_2
Xtap_48_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[5\].RFW.BIT\[29\].FF REGF\[5\].RFW.CG\[3\]/GCLK DW[29] VGND VGND VPWR VPWR
+ REGF\[5\].RFW.BIT\[29\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[11\].RFW.BIT\[19\].FF REGF\[11\].RFW.CG\[2\]/GCLK DW[19] VGND VGND VPWR VPWR
+ REGF\[11\].RFW.BIT\[19\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[1\].RFW.BIT\[31\].FF REGF\[1\].RFW.CG\[3\]/GCLK DW[31] VGND VGND VPWR VPWR
+ REGF\[1\].RFW.BIT\[31\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_12_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[17\].RFW.BIT\[13\].FF REGF\[17\].RFW.CG\[1\]/GCLK DW[13] VGND VGND VPWR VPWR
+ REGF\[17\].RFW.BIT\[13\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[11\].RFW.CG\[1\] CLK REGF\[11\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[11\].RFW.CG\[1\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[7\].RFW.BIT\[2\].OBUF2 REGF\[7\].RFW.BIT\[2\].FF/Q REGF\[7\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[2] sky130_fd_sc_hd__ebufn_2
Xfill_36_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_36_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDEC2.D2.AND5 DEC2.D2.AND7/B DEC2.D2.AND7/A DEC2.D2.AND7/C DEC2.D2.AND7/D VGND VGND
+ VPWR VPWR DEC2.D2.AND5/X sky130_fd_sc_hd__and4b_2
Xfill_52_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_52_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[10\].RFW.BIT\[1\].OBUF2 REGF\[10\].RFW.BIT\[1\].FF/Q REGF\[10\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[1] sky130_fd_sc_hd__ebufn_2
Xfill_8_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[19\].RFW.BIT\[28\].OBUF1 REGF\[19\].RFW.BIT\[28\].FF/Q REGF\[19\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[28] sky130_fd_sc_hd__ebufn_2
Xfill_8_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_8_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[28\].RFW.BIT\[8\].OBUF1 REGF\[28\].RFW.BIT\[8\].FF/Q REGF\[28\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[8] sky130_fd_sc_hd__ebufn_2
XREGF\[22\].RFW.BIT\[29\].FF REGF\[22\].RFW.CG\[3\]/GCLK DW[29] VGND VGND VPWR VPWR
+ REGF\[22\].RFW.BIT\[29\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[24\].RFW.BIT\[17\].OBUF1 REGF\[24\].RFW.BIT\[17\].FF/Q REGF\[24\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[17] sky130_fd_sc_hd__ebufn_2
XREGF\[25\].RFW.BIT\[30\].OBUF1 REGF\[25\].RFW.BIT\[30\].FF/Q REGF\[25\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[30] sky130_fd_sc_hd__ebufn_2
Xfill_40_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[28\].RFW.BIT\[23\].FF REGF\[28\].RFW.CG\[2\]/GCLK DW[23] VGND VGND VPWR VPWR
+ REGF\[28\].RFW.BIT\[23\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_33_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_26_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfill_19_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[19\].RFW.BIT\[3\].OBUF2 REGF\[19\].RFW.BIT\[3\].FF/Q REGF\[19\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[3] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.BIT\[6\].OBUF1 REGF\[21\].RFW.BIT\[6\].FF/Q REGF\[21\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[6] sky130_fd_sc_hd__ebufn_2
Xtap_48_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC1.D1.ENBUF DEC1.D.AND1/X VGND VGND VPWR VPWR DEC1.D1.AND7/D sky130_fd_sc_hd__clkbuf_2
XREGF\[9\].RFW.BIT\[2\].OBUF2 REGF\[9\].RFW.BIT\[2\].FF/Q REGF\[9\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[2] sky130_fd_sc_hd__ebufn_2
Xtap_18_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_57_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[2\].RFW.BIT\[14\].FF REGF\[2\].RFW.CG\[1\]/GCLK DW[14] VGND VGND VPWR VPWR
+ REGF\[2\].RFW.BIT\[14\].FF/Q sky130_fd_sc_hd__dfxtp_1
XDEC1.D3.AND7 DEC1.D3.AND7/A DEC1.D3.AND7/B DEC1.D3.AND7/C DEC1.D3.AND7/D VGND VGND
+ VPWR VPWR DEC1.D3.AND7/X sky130_fd_sc_hd__and4_2
XREGF\[28\].RFW.BIT\[18\].OBUF2 REGF\[28\].RFW.BIT\[18\].FF/Q REGF\[28\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[18] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.BIT\[31\].OBUF2 REGF\[29\].RFW.BIT\[31\].FF/Q REGF\[29\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[31] sky130_fd_sc_hd__ebufn_2
Xtap_34_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.BIT\[1\].OBUF2 REGF\[12\].RFW.BIT\[1\].FF/Q REGF\[12\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[1] sky130_fd_sc_hd__ebufn_2
Xtap_50_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.BIT\[23\].OBUF1 REGF\[6\].RFW.BIT\[23\].FF/Q REGF\[6\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[23] sky130_fd_sc_hd__ebufn_2
Xfill_22_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_22_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_22_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.BIT\[16\].OBUF1 REGF\[18\].RFW.BIT\[16\].FF/Q REGF\[18\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[16] sky130_fd_sc_hd__ebufn_2
XREGF\[2\].RFW.BIT\[0\].OBUF2 REGF\[2\].RFW.BIT\[0\].FF/Q REGF\[2\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[0] sky130_fd_sc_hd__ebufn_2
Xfill_47_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_47_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_47_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_47_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_12_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[23\].RFW.BIT\[6\].OBUF1 REGF\[23\].RFW.BIT\[6\].FF/Q REGF\[23\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[6] sky130_fd_sc_hd__ebufn_2
XREGF\[30\].RFW.BIT\[23\].OBUF2 REGF\[30\].RFW.BIT\[23\].FF/Q REGF\[30\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[23] sky130_fd_sc_hd__ebufn_2
XREGF\[14\].RFW.BIT\[1\].OBUF2 REGF\[14\].RFW.BIT\[1\].FF/Q REGF\[14\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[1] sky130_fd_sc_hd__ebufn_2
XREGF\[2\].RFW.BIT\[26\].OBUF1 REGF\[2\].RFW.BIT\[26\].FF/Q REGF\[2\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[26] sky130_fd_sc_hd__ebufn_2
XREGF\[14\].RFW.BIT\[19\].OBUF1 REGF\[14\].RFW.BIT\[19\].FF/Q REGF\[14\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[19] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.BIT\[19\].FF REGF\[18\].RFW.CG\[2\]/GCLK DW[19] VGND VGND VPWR VPWR
+ REGF\[18\].RFW.BIT\[19\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[8\].RFW.BIT\[31\].FF REGF\[8\].RFW.CG\[3\]/GCLK DW[31] VGND VGND VPWR VPWR
+ REGF\[8\].RFW.BIT\[31\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[14\].RFW.BIT\[21\].FF REGF\[14\].RFW.CG\[2\]/GCLK DW[21] VGND VGND VPWR VPWR
+ REGF\[14\].RFW.BIT\[21\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_31_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[30\].RFW.BIT\[24\].FF REGF\[30\].RFW.CG\[3\]/GCLK DW[24] VGND VGND VPWR VPWR
+ REGF\[30\].RFW.BIT\[24\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[20\].RFW.BIT\[21\].OBUF1 REGF\[20\].RFW.BIT\[21\].FF/Q REGF\[20\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[21] sky130_fd_sc_hd__ebufn_2
XREGF\[6\].RFW.INV1\[2\] DEC0.D0.AND6/X VGND VGND VPWR VPWR REGF\[6\].RFW.INV1\[2\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[4\].RFW.BIT\[0\].OBUF2 REGF\[4\].RFW.BIT\[0\].FF/Q REGF\[4\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[0] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[11\].OBUF1 REGF\[5\].RFW.BIT\[11\].FF/Q REGF\[5\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[11] sky130_fd_sc_hd__ebufn_2
Xtap_60_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_46_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.BIT\[27\].OBUF2 REGF\[6\].RFW.BIT\[27\].FF/Q REGF\[6\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[27] sky130_fd_sc_hd__ebufn_2
XREGF\[25\].RFW.BIT\[6\].OBUF1 REGF\[25\].RFW.BIT\[6\].FF/Q REGF\[25\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[6] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.INV1\[0\] DEC0.D3.AND2/X VGND VGND VPWR VPWR REGF\[26\].RFW.INV1\[0\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[29\].RFW.BIT\[29\].FF REGF\[29\].RFW.CG\[3\]/GCLK DW[29] VGND VGND VPWR VPWR
+ REGF\[29\].RFW.BIT\[29\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[25\].RFW.BIT\[31\].FF REGF\[25\].RFW.CG\[3\]/GCLK DW[31] VGND VGND VPWR VPWR
+ REGF\[25\].RFW.BIT\[31\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_17_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_17_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_17_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_17_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_17_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[24\].RFW.BIT\[22\].OBUF2 REGF\[24\].RFW.BIT\[22\].FF/Q REGF\[24\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[22] sky130_fd_sc_hd__ebufn_2
Xfill_33_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_33_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[16\].RFW.BIT\[1\].OBUF2 REGF\[16\].RFW.BIT\[1\].FF/Q REGF\[16\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[1] sky130_fd_sc_hd__ebufn_2
Xfill_33_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_33_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[9\].RFW.BIT\[12\].OBUF2 REGF\[9\].RFW.BIT\[12\].FF/Q REGF\[9\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[12] sky130_fd_sc_hd__ebufn_2
XREGF\[1\].RFW.BIT\[14\].OBUF1 REGF\[1\].RFW.BIT\[14\].FF/Q REGF\[1\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[14] sky130_fd_sc_hd__ebufn_2
Xfill_58_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[14\].RFW.BIT\[20\].OBUF1 REGF\[14\].RFW.BIT\[20\].FF/Q REGF\[14\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[20] sky130_fd_sc_hd__ebufn_2
Xfill_5_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_5_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_5_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_5_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[15\].RFW.BIT\[1\].FF REGF\[15\].RFW.CG\[0\]/GCLK DW[1] VGND VGND VPWR VPWR
+ REGF\[15\].RFW.BIT\[1\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[6\].RFW.BIT\[0\].OBUF2 REGF\[6\].RFW.BIT\[0\].FF/Q REGF\[6\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[0] sky130_fd_sc_hd__ebufn_2
XREGF\[9\].RFW.BIT\[14\].FF REGF\[9\].RFW.CG\[1\]/GCLK DW[14] VGND VGND VPWR VPWR
+ REGF\[9\].RFW.BIT\[14\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_10_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_8_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[25\].OBUF2 REGF\[20\].RFW.BIT\[25\].FF/Q REGF\[20\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[25] sky130_fd_sc_hd__ebufn_2
XREGF\[14\].RFW.BIT\[3\].FF REGF\[14\].RFW.CG\[0\]/GCLK DW[3] VGND VGND VPWR VPWR
+ REGF\[14\].RFW.BIT\[3\].FF/Q sky130_fd_sc_hd__dfxtp_1
XDEC0.D.AND3 RA[4] RA[3] DEC0.TIE/HI VGND VGND VPWR VPWR DEC0.D.AND3/X sky130_fd_sc_hd__and3_4
XREGF\[27\].RFW.BIT\[6\].OBUF1 REGF\[27\].RFW.BIT\[6\].FF/Q REGF\[27\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[6] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[15\].OBUF2 REGF\[5\].RFW.BIT\[15\].FF/Q REGF\[5\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[15] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.BIT\[21\].OBUF2 REGF\[18\].RFW.BIT\[21\].FF/Q REGF\[18\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[21] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.BIT\[1\].OBUF2 REGF\[18\].RFW.BIT\[1\].FF/Q REGF\[18\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[1] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[14\].FF REGF\[26\].RFW.CG\[1\]/GCLK DW[14] VGND VGND VPWR VPWR
+ REGF\[26\].RFW.BIT\[14\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[10\].RFW.BIT\[23\].OBUF1 REGF\[10\].RFW.BIT\[23\].FF/Q REGF\[10\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[23] sky130_fd_sc_hd__ebufn_2
XREGF\[23\].RFW.BIT\[10\].OBUF2 REGF\[23\].RFW.BIT\[10\].FF/Q REGF\[23\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[10] sky130_fd_sc_hd__ebufn_2
XREGF\[13\].RFW.BIT\[5\].FF REGF\[13\].RFW.CG\[0\]/GCLK DW[5] VGND VGND VPWR VPWR
+ REGF\[13\].RFW.BIT\[5\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[20\].RFW.BIT\[4\].OBUF1 REGF\[20\].RFW.BIT\[4\].FF/Q REGF\[20\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[4] sky130_fd_sc_hd__ebufn_2
XREGF\[8\].RFW.CGAND DEC2.D1.AND0/Y WE VGND VGND VPWR VPWR REGF\[8\].RFW.CGAND/X sky130_fd_sc_hd__and2_1
Xtap_44_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[8\].RFW.BIT\[0\].OBUF2 REGF\[8\].RFW.BIT\[0\].FF/Q REGF\[8\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[0] sky130_fd_sc_hd__ebufn_2
Xtap_37_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.CG\[0\] CLK REGF\[31\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[31\].RFW.CG\[0\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_56_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[28\].RFW.BIT\[1\].FF REGF\[28\].RFW.CG\[0\]/GCLK DW[1] VGND VGND VPWR VPWR
+ REGF\[28\].RFW.BIT\[1\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[15\].RFW.BIT\[27\].FF REGF\[15\].RFW.CG\[3\]/GCLK DW[27] VGND VGND VPWR VPWR
+ REGF\[15\].RFW.BIT\[27\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[12\].RFW.BIT\[7\].FF REGF\[12\].RFW.CG\[0\]/GCLK DW[7] VGND VGND VPWR VPWR
+ REGF\[12\].RFW.BIT\[7\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_28_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_28_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_28_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.INV2\[1\] DEC1.D2.AND4/X VGND VGND VPWR VPWR REGF\[20\].RFW.INV2\[1\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[1\].RFW.BIT\[18\].OBUF2 REGF\[1\].RFW.BIT\[18\].FF/Q REGF\[1\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[18] sky130_fd_sc_hd__ebufn_2
Xfill_44_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[2\].RFW.BIT\[31\].OBUF2 REGF\[2\].RFW.BIT\[31\].FF/Q REGF\[2\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[31] sky130_fd_sc_hd__ebufn_2
Xfill_44_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[29\].RFW.BIT\[6\].OBUF1 REGF\[29\].RFW.BIT\[6\].FF/Q REGF\[29\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[6] sky130_fd_sc_hd__ebufn_2
XREGF\[14\].RFW.BIT\[24\].OBUF2 REGF\[14\].RFW.BIT\[24\].FF/Q REGF\[14\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[24] sky130_fd_sc_hd__ebufn_2
Xfill_60_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_60_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[27\].RFW.BIT\[3\].FF REGF\[27\].RFW.CG\[0\]/GCLK DW[3] VGND VGND VPWR VPWR
+ REGF\[27\].RFW.BIT\[3\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[11\].RFW.BIT\[9\].FF REGF\[11\].RFW.CG\[1\]/GCLK DW[9] VGND VGND VPWR VPWR
+ REGF\[11\].RFW.BIT\[9\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_58_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[9\].RFW.CG\[3\] CLK REGF\[9\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[9\].RFW.CG\[3\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[20\].RFW.CG\[3\] CLK REGF\[20\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[20\].RFW.CG\[3\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_6_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[22\].RFW.BIT\[4\].OBUF1 REGF\[22\].RFW.BIT\[4\].FF/Q REGF\[22\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[4] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[5\].FF REGF\[26\].RFW.CG\[0\]/GCLK DW[5] VGND VGND VPWR VPWR
+ REGF\[26\].RFW.BIT\[5\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[10\].RFW.BIT\[27\].OBUF2 REGF\[10\].RFW.BIT\[27\].FF/Q REGF\[10\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[27] sky130_fd_sc_hd__ebufn_2
Xtap_30_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[25\].RFW.BIT\[7\].FF REGF\[25\].RFW.CG\[0\]/GCLK DW[7] VGND VGND VPWR VPWR
+ REGF\[25\].RFW.BIT\[7\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_26_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[8\].OBUF2 REGF\[20\].RFW.BIT\[8\].FF/Q REGF\[20\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[8] sky130_fd_sc_hd__ebufn_2
XREGF\[6\].RFW.BIT\[22\].FF REGF\[6\].RFW.CG\[2\]/GCLK DW[22] VGND VGND VPWR VPWR
+ REGF\[6\].RFW.BIT\[22\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[12\].RFW.BIT\[12\].FF REGF\[12\].RFW.CG\[1\]/GCLK DW[12] VGND VGND VPWR VPWR
+ REGF\[12\].RFW.BIT\[12\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_42_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[8\].RFW.CG\[0\] CLK REGF\[8\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[8\].RFW.CG\[0\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[13\].RFW.BIT\[12\].OBUF2 REGF\[13\].RFW.BIT\[12\].FF/Q REGF\[13\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[12] sky130_fd_sc_hd__ebufn_2
Xfill_14_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_14_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_14_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_30_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_30_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_30_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[24\].RFW.BIT\[9\].FF REGF\[24\].RFW.CG\[1\]/GCLK DW[9] VGND VGND VPWR VPWR
+ REGF\[24\].RFW.BIT\[9\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[31\].RFW.BIT\[26\].OBUF1 REGF\[31\].RFW.BIT\[26\].FF/Q REGF\[31\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[26] sky130_fd_sc_hd__ebufn_2
XDEC0.D0.AND1 DEC0.D0.AND7/C DEC0.D0.AND7/B DEC0.D0.AND7/A DEC0.D0.AND7/D VGND VGND
+ VPWR VPWR DEC0.D0.AND1/X sky130_fd_sc_hd__and4bb_2
Xtap_42_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[15\].RFW.INV2\[2\] DEC1.D1.AND7/X VGND VGND VPWR VPWR REGF\[15\].RFW.INV2\[2\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[24\].RFW.BIT\[4\].OBUF1 REGF\[24\].RFW.BIT\[4\].FF/Q REGF\[24\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[4] sky130_fd_sc_hd__ebufn_2
Xfill_39_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[29\].RFW.BIT\[22\].OBUF1 REGF\[29\].RFW.BIT\[22\].FF/Q REGF\[29\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[22] sky130_fd_sc_hd__ebufn_2
Xfill_55_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_2_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_55_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_55_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_55_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_2_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_2_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[18\].RFW.CGAND DEC2.D2.AND2/X WE VGND VGND VPWR VPWR REGF\[18\].RFW.CGAND/X
+ sky130_fd_sc_hd__and2_1
XREGF\[23\].RFW.BIT\[22\].FF REGF\[23\].RFW.CG\[2\]/GCLK DW[22] VGND VGND VPWR VPWR
+ REGF\[23\].RFW.BIT\[22\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[22\].RFW.BIT\[8\].OBUF2 REGF\[22\].RFW.BIT\[8\].FF/Q REGF\[22\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[8] sky130_fd_sc_hd__ebufn_2
XREGF\[9\].RFW.BIT\[6\].FF REGF\[9\].RFW.CG\[0\]/GCLK DW[6] VGND VGND VPWR VPWR REGF\[9\].RFW.BIT\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xfill_56_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_49_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDEC2.D3.ABUF\[2\] RW[2] VGND VGND VPWR VPWR DEC2.D3.AND7/C sky130_fd_sc_hd__clkbuf_2
Xfill_4_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[25\].RFW.BIT\[25\].OBUF1 REGF\[25\].RFW.BIT\[25\].FF/Q REGF\[25\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[25] sky130_fd_sc_hd__ebufn_2
XREGF\[8\].RFW.BIT\[8\].FF REGF\[8\].RFW.CG\[1\]/GCLK DW[8] VGND VGND VPWR VPWR REGF\[8\].RFW.BIT\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[30\].RFW.BIT\[14\].OBUF1 REGF\[30\].RFW.BIT\[14\].FF/Q REGF\[30\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[14] sky130_fd_sc_hd__ebufn_2
XREGF\[11\].RFW.INV1\[3\] DEC0.D1.AND3/X VGND VGND VPWR VPWR REGF\[11\].RFW.INV1\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[26\].RFW.BIT\[4\].OBUF1 REGF\[26\].RFW.BIT\[4\].FF/Q REGF\[26\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[4] sky130_fd_sc_hd__ebufn_2
Xtap_21_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_14_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[28\].RFW.BIT\[10\].OBUF1 REGF\[28\].RFW.BIT\[10\].FF/Q REGF\[28\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[10] sky130_fd_sc_hd__ebufn_2
Xtap_7_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgenblk1.RFW0.BIT\[3\].OBUF2 genblk1.RFW0.TIE\[4\]/LO genblk1.RFW0.INV2\[0\]/Y VGND
+ VGND VPWR VPWR DB[3] sky130_fd_sc_hd__ebufn_2
Xfill_25_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_25_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_25_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_25_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[24\].RFW.BIT\[8\].OBUF2 REGF\[24\].RFW.BIT\[8\].FF/Q REGF\[24\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[8] sky130_fd_sc_hd__ebufn_2
Xfill_41_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_41_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_41_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[29\].RFW.BIT\[26\].OBUF2 REGF\[29\].RFW.BIT\[26\].FF/Q REGF\[29\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[26] sky130_fd_sc_hd__ebufn_2
Xfill_41_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_41_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_41_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[21\].RFW.BIT\[28\].OBUF1 REGF\[21\].RFW.BIT\[28\].FF/Q REGF\[21\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[28] sky130_fd_sc_hd__ebufn_2
XREGF\[7\].RFW.BIT\[31\].OBUF1 REGF\[7\].RFW.BIT\[31\].FF/Q REGF\[7\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[31] sky130_fd_sc_hd__ebufn_2
XREGF\[6\].RFW.BIT\[18\].OBUF1 REGF\[6\].RFW.BIT\[18\].FF/Q REGF\[6\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[18] sky130_fd_sc_hd__ebufn_2
Xfill_42_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[7\].RFW.BIT\[28\].FF REGF\[7\].RFW.CG\[3\]/GCLK DW[28] VGND VGND VPWR VPWR
+ REGF\[7\].RFW.BIT\[28\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[13\].RFW.BIT\[18\].FF REGF\[13\].RFW.CG\[2\]/GCLK DW[18] VGND VGND VPWR VPWR
+ REGF\[13\].RFW.BIT\[18\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[19\].RFW.BIT\[24\].OBUF1 REGF\[19\].RFW.BIT\[24\].FF/Q REGF\[19\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[24] sky130_fd_sc_hd__ebufn_2
Xfill_28_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[28\].RFW.BIT\[4\].OBUF1 REGF\[28\].RFW.BIT\[4\].FF/Q REGF\[28\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[4] sky130_fd_sc_hd__ebufn_2
XREGF\[3\].RFW.BIT\[30\].FF REGF\[3\].RFW.CG\[3\]/GCLK DW[30] VGND VGND VPWR VPWR
+ REGF\[3\].RFW.BIT\[30\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[24\].RFW.BIT\[13\].OBUF1 REGF\[24\].RFW.BIT\[13\].FF/Q REGF\[24\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[13] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.BIT\[12\].FF REGF\[19\].RFW.CG\[1\]/GCLK DW[12] VGND VGND VPWR VPWR
+ REGF\[19\].RFW.BIT\[12\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_61_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[25\].RFW.BIT\[29\].OBUF2 REGF\[25\].RFW.BIT\[29\].FF/Q REGF\[25\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[29] sky130_fd_sc_hd__ebufn_2
XREGF\[2\].RFW.INV2\[0\] DEC1.D0.AND2/X VGND VGND VPWR VPWR REGF\[2\].RFW.INV2\[0\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[26\].RFW.BIT\[8\].OBUF2 REGF\[26\].RFW.BIT\[8\].FF/Q REGF\[26\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[8] sky130_fd_sc_hd__ebufn_2
XREGF\[30\].RFW.BIT\[18\].OBUF2 REGF\[30\].RFW.BIT\[18\].FF/Q REGF\[30\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[18] sky130_fd_sc_hd__ebufn_2
XREGF\[31\].RFW.BIT\[31\].OBUF2 REGF\[31\].RFW.BIT\[31\].FF/Q REGF\[31\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[31] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.BIT\[2\].OBUF1 REGF\[21\].RFW.BIT\[2\].FF/Q REGF\[21\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[2] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[28\].FF REGF\[24\].RFW.CG\[3\]/GCLK DW[28] VGND VGND VPWR VPWR
+ REGF\[24\].RFW.BIT\[28\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[20\].RFW.BIT\[30\].FF REGF\[20\].RFW.CG\[3\]/GCLK DW[30] VGND VGND VPWR VPWR
+ REGF\[20\].RFW.BIT\[30\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[15\].RFW.BIT\[27\].OBUF1 REGF\[15\].RFW.BIT\[27\].FF/Q REGF\[15\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[27] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.BIT\[14\].OBUF2 REGF\[28\].RFW.BIT\[14\].FF/Q REGF\[28\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[14] sky130_fd_sc_hd__ebufn_2
Xfill_11_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_11_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[16\].OBUF1 REGF\[20\].RFW.BIT\[16\].FF/Q REGF\[20\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[16] sky130_fd_sc_hd__ebufn_2
Xfill_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_11_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_11_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_48_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.BIT\[12\].OBUF1 REGF\[18\].RFW.BIT\[12\].FF/Q REGF\[18\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[12] sky130_fd_sc_hd__ebufn_2
Xfill_36_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_36_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_36_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[4\].RFW.BIT\[13\].FF REGF\[4\].RFW.CG\[1\]/GCLK DW[13] VGND VGND VPWR VPWR
+ REGF\[4\].RFW.BIT\[13\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_52_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_52_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC2.D2.AND6 DEC2.D2.AND7/A DEC2.D2.AND7/B DEC2.D2.AND7/C DEC2.D2.AND7/D VGND VGND
+ VPWR VPWR DEC2.D2.AND6/X sky130_fd_sc_hd__and4b_2
Xfill_8_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_8_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_8_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[19\].RFW.BIT\[28\].OBUF2 REGF\[19\].RFW.BIT\[28\].FF/Q REGF\[19\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[28] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.BIT\[8\].OBUF2 REGF\[28\].RFW.BIT\[8\].FF/Q REGF\[28\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[8] sky130_fd_sc_hd__ebufn_2
XREGF\[23\].RFW.BIT\[2\].OBUF1 REGF\[23\].RFW.BIT\[2\].FF/Q REGF\[23\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[2] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[17\].OBUF2 REGF\[24\].RFW.BIT\[17\].FF/Q REGF\[24\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[17] sky130_fd_sc_hd__ebufn_2
XREGF\[25\].RFW.BIT\[30\].OBUF2 REGF\[25\].RFW.BIT\[30\].FF/Q REGF\[25\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[30] sky130_fd_sc_hd__ebufn_2
Xfill_40_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_33_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_26_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_19_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XREGF\[2\].RFW.BIT\[22\].OBUF1 REGF\[2\].RFW.BIT\[22\].FF/Q REGF\[2\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[22] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.BIT\[13\].FF REGF\[21\].RFW.CG\[1\]/GCLK DW[13] VGND VGND VPWR VPWR
+ REGF\[21\].RFW.BIT\[13\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[14\].RFW.BIT\[15\].OBUF1 REGF\[14\].RFW.BIT\[15\].FF/Q REGF\[14\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[15] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.BIT\[6\].OBUF2 REGF\[21\].RFW.BIT\[6\].FF/Q REGF\[21\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[6] sky130_fd_sc_hd__ebufn_2
XREGF\[10\].RFW.BIT\[26\].FF REGF\[10\].RFW.CG\[3\]/GCLK DW[26] VGND VGND VPWR VPWR
+ REGF\[10\].RFW.BIT\[26\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[16\].RFW.BIT\[20\].FF REGF\[16\].RFW.CG\[2\]/GCLK DW[20] VGND VGND VPWR VPWR
+ REGF\[16\].RFW.BIT\[20\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_50_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.BIT\[23\].OBUF2 REGF\[6\].RFW.BIT\[23\].FF/Q REGF\[6\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[23] sky130_fd_sc_hd__ebufn_2
XREGF\[22\].RFW.BIT\[0\].FF REGF\[22\].RFW.CG\[0\]/GCLK DW[0] VGND VGND VPWR VPWR
+ REGF\[22\].RFW.BIT\[0\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_22_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_22_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_22_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[25\].RFW.BIT\[2\].OBUF1 REGF\[25\].RFW.BIT\[2\].FF/Q REGF\[25\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[2] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.BIT\[16\].OBUF2 REGF\[18\].RFW.BIT\[16\].FF/Q REGF\[18\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[16] sky130_fd_sc_hd__ebufn_2
XREGF\[11\].RFW.BIT\[31\].OBUF1 REGF\[11\].RFW.BIT\[31\].FF/Q REGF\[11\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[31] sky130_fd_sc_hd__ebufn_2
XREGF\[10\].RFW.BIT\[18\].OBUF1 REGF\[10\].RFW.BIT\[18\].FF/Q REGF\[10\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[18] sky130_fd_sc_hd__ebufn_2
Xfill_47_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_47_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_47_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_47_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_47_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[21\].RFW.BIT\[2\].FF REGF\[21\].RFW.CG\[0\]/GCLK DW[2] VGND VGND VPWR VPWR
+ REGF\[21\].RFW.BIT\[2\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[1\].RFW.BIT\[10\].OBUF1 REGF\[1\].RFW.BIT\[10\].FF/Q REGF\[1\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[10] sky130_fd_sc_hd__ebufn_2
Xfill_12_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[23\].RFW.BIT\[6\].OBUF2 REGF\[23\].RFW.BIT\[6\].FF/Q REGF\[23\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[6] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[30\].FF REGF\[27\].RFW.CG\[3\]/GCLK DW[30] VGND VGND VPWR VPWR
+ REGF\[27\].RFW.BIT\[30\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[9\].RFW.INV1\[3\] DEC0.D1.AND1/X VGND VGND VPWR VPWR REGF\[9\].RFW.INV1\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[2\].RFW.BIT\[26\].OBUF2 REGF\[2\].RFW.BIT\[26\].FF/Q REGF\[2\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[26] sky130_fd_sc_hd__ebufn_2
XREGF\[20\].RFW.BIT\[4\].FF REGF\[20\].RFW.CG\[0\]/GCLK DW[4] VGND VGND VPWR VPWR
+ REGF\[20\].RFW.BIT\[4\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[14\].RFW.BIT\[19\].OBUF2 REGF\[14\].RFW.BIT\[19\].FF/Q REGF\[14\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[19] sky130_fd_sc_hd__ebufn_2
Xfill_31_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[20\].RFW.BIT\[21\].OBUF2 REGF\[20\].RFW.BIT\[21\].FF/Q REGF\[20\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[21] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[2\].OBUF1 REGF\[27\].RFW.BIT\[2\].FF/Q REGF\[27\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[2] sky130_fd_sc_hd__ebufn_2
Xfill_24_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[5\].RFW.BIT\[19\].FF REGF\[5\].RFW.CG\[2\]/GCLK DW[19] VGND VGND VPWR VPWR
+ REGF\[5\].RFW.BIT\[19\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[13\].RFW.INV1\[0\] DEC0.D1.AND5/X VGND VGND VPWR VPWR REGF\[13\].RFW.INV1\[0\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[5\].RFW.BIT\[11\].OBUF2 REGF\[5\].RFW.BIT\[11\].FF/Q REGF\[5\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[11] sky130_fd_sc_hd__ebufn_2
XREGF\[1\].RFW.BIT\[21\].FF REGF\[1\].RFW.CG\[2\]/GCLK DW[21] VGND VGND VPWR VPWR
+ REGF\[1\].RFW.BIT\[21\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_60_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[7\].RFW.CGAND DEC2.D0.AND7/X WE VGND VGND VPWR VPWR REGF\[7\].RFW.CGAND/X sky130_fd_sc_hd__and2_1
XREGF\[29\].RFW.INV1\[1\] DEC0.D3.AND5/X VGND VGND VPWR VPWR REGF\[29\].RFW.INV1\[1\]/Y
+ sky130_fd_sc_hd__inv_4
Xtap_46_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[25\].RFW.BIT\[6\].OBUF2 REGF\[25\].RFW.BIT\[6\].FF/Q REGF\[25\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[6] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[1\].FF REGF\[5\].RFW.CG\[0\]/GCLK DW[1] VGND VGND VPWR VPWR REGF\[5\].RFW.BIT\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[20\].RFW.BIT\[0\].OBUF1 REGF\[20\].RFW.BIT\[0\].FF/Q REGF\[20\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[0] sky130_fd_sc_hd__ebufn_2
Xfill_17_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_17_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_17_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_17_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_17_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[22\].RFW.BIT\[19\].FF REGF\[22\].RFW.CG\[2\]/GCLK DW[19] VGND VGND VPWR VPWR
+ REGF\[22\].RFW.BIT\[19\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_33_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_33_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_33_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_33_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[28\].RFW.BIT\[13\].FF REGF\[28\].RFW.CG\[1\]/GCLK DW[13] VGND VGND VPWR VPWR
+ REGF\[28\].RFW.BIT\[13\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[1\].RFW.BIT\[14\].OBUF2 REGF\[1\].RFW.BIT\[14\].FF/Q REGF\[1\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[14] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.BIT\[3\].FF REGF\[4\].RFW.CG\[0\]/GCLK DW[3] VGND VGND VPWR VPWR REGF\[4\].RFW.BIT\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[29\].RFW.BIT\[2\].OBUF1 REGF\[29\].RFW.BIT\[2\].FF/Q REGF\[29\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[2] sky130_fd_sc_hd__ebufn_2
Xfill_58_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_58_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[14\].RFW.BIT\[20\].OBUF2 REGF\[14\].RFW.BIT\[20\].FF/Q REGF\[14\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[20] sky130_fd_sc_hd__ebufn_2
Xfill_5_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_5_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_5_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_5_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_5_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[5\].RFW.CG\[2\] CLK REGF\[5\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[5\].RFW.CG\[2\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_10_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_8_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC1.D0.ENBUF DEC1.D.AND0/Y VGND VGND VPWR VPWR DEC1.D0.AND7/D sky130_fd_sc_hd__clkbuf_2
XREGF\[17\].RFW.BIT\[26\].FF REGF\[17\].RFW.CG\[3\]/GCLK DW[26] VGND VGND VPWR VPWR
+ REGF\[17\].RFW.BIT\[26\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[3\].RFW.BIT\[5\].FF REGF\[3\].RFW.CG\[0\]/GCLK DW[5] VGND VGND VPWR VPWR REGF\[3\].RFW.BIT\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[29\].RFW.BIT\[17\].OBUF1 REGF\[29\].RFW.BIT\[17\].FF/Q REGF\[29\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[17] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[6\].OBUF2 REGF\[27\].RFW.BIT\[6\].FF/Q REGF\[27\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[6] sky130_fd_sc_hd__ebufn_2
XREGF\[22\].RFW.BIT\[0\].OBUF1 REGF\[22\].RFW.BIT\[0\].FF/Q REGF\[22\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[0] sky130_fd_sc_hd__ebufn_2
XREGF\[2\].RFW.BIT\[7\].FF REGF\[2\].RFW.CG\[0\]/GCLK DW[7] VGND VGND VPWR VPWR REGF\[2\].RFW.BIT\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[31\].RFW.BIT\[8\].FF REGF\[31\].RFW.CG\[1\]/GCLK DW[8] VGND VGND VPWR VPWR
+ REGF\[31\].RFW.BIT\[8\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[10\].RFW.BIT\[23\].OBUF2 REGF\[10\].RFW.BIT\[23\].FF/Q REGF\[10\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[23] sky130_fd_sc_hd__ebufn_2
XREGF\[20\].RFW.BIT\[4\].OBUF2 REGF\[20\].RFW.BIT\[4\].FF/Q REGF\[20\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[4] sky130_fd_sc_hd__ebufn_2
XREGF\[23\].RFW.INV2\[2\] DEC1.D2.AND7/X VGND VGND VPWR VPWR REGF\[23\].RFW.INV2\[2\]/Y
+ sky130_fd_sc_hd__inv_4
Xtap_44_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_37_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[1\].RFW.BIT\[9\].FF REGF\[1\].RFW.CG\[1\]/GCLK DW[9] VGND VGND VPWR VPWR REGF\[1\].RFW.BIT\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xtap_56_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_28_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_28_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_28_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.BIT\[22\].OBUF1 REGF\[31\].RFW.BIT\[22\].FF/Q REGF\[31\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[22] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.CGAND DEC2.D2.AND1/X WE VGND VGND VPWR VPWR REGF\[17\].RFW.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_44_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_44_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_44_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[2\].RFW.BIT\[27\].FF REGF\[2\].RFW.CG\[3\]/GCLK DW[27] VGND VGND VPWR VPWR
+ REGF\[2\].RFW.BIT\[27\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[24\].RFW.BIT\[0\].OBUF1 REGF\[24\].RFW.BIT\[0\].FF/Q REGF\[24\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[0] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.BIT\[6\].OBUF2 REGF\[29\].RFW.BIT\[6\].FF/Q REGF\[29\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[6] sky130_fd_sc_hd__ebufn_2
Xfill_60_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_60_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[8\].RFW.BIT\[21\].FF REGF\[8\].RFW.CG\[2\]/GCLK DW[21] VGND VGND VPWR VPWR
+ REGF\[8\].RFW.BIT\[21\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[14\].RFW.BIT\[11\].FF REGF\[14\].RFW.CG\[1\]/GCLK DW[11] VGND VGND VPWR VPWR
+ REGF\[14\].RFW.BIT\[11\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[30\].RFW.BIT\[14\].FF REGF\[30\].RFW.CG\[1\]/GCLK DW[14] VGND VGND VPWR VPWR
+ REGF\[30\].RFW.BIT\[14\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[31\].RFW.BIT\[9\].OBUF1 REGF\[31\].RFW.BIT\[9\].FF/Q REGF\[31\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[9] sky130_fd_sc_hd__ebufn_2
Xfill_58_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_6_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[22\].RFW.BIT\[4\].OBUF2 REGF\[22\].RFW.BIT\[4\].FF/Q REGF\[22\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[4] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.CG\[1\] CLK REGF\[19\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[19\].RFW.CG\[1\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[29\].RFW.BIT\[19\].FF REGF\[29\].RFW.CG\[2\]/GCLK DW[19] VGND VGND VPWR VPWR
+ REGF\[29\].RFW.BIT\[19\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[7\].RFW.BIT\[26\].OBUF1 REGF\[7\].RFW.BIT\[26\].FF/Q REGF\[7\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[26] sky130_fd_sc_hd__ebufn_2
XREGF\[25\].RFW.BIT\[21\].FF REGF\[25\].RFW.CG\[2\]/GCLK DW[21] VGND VGND VPWR VPWR
+ REGF\[25\].RFW.BIT\[21\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[19\].RFW.BIT\[19\].OBUF1 REGF\[19\].RFW.BIT\[19\].FF/Q REGF\[19\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[19] sky130_fd_sc_hd__ebufn_2
XREGF\[25\].RFW.BIT\[21\].OBUF1 REGF\[25\].RFW.BIT\[21\].FF/Q REGF\[25\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[21] sky130_fd_sc_hd__ebufn_2
Xtap_16_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[26\].RFW.BIT\[0\].OBUF1 REGF\[26\].RFW.BIT\[0\].FF/Q REGF\[26\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[0] sky130_fd_sc_hd__ebufn_2
XREGF\[30\].RFW.BIT\[10\].OBUF1 REGF\[30\].RFW.BIT\[10\].FF/Q REGF\[30\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[10] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.INV2\[3\] DEC1.D2.AND2/X VGND VGND VPWR VPWR REGF\[18\].RFW.INV2\[3\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_14_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_14_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_14_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_30_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_30_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[31\].RFW.BIT\[26\].OBUF2 REGF\[31\].RFW.BIT\[26\].FF/Q REGF\[31\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[26] sky130_fd_sc_hd__ebufn_2
XDEC0.D0.AND2 DEC0.D0.AND7/C DEC0.D0.AND7/A DEC0.D0.AND7/B DEC0.D0.AND7/D VGND VGND
+ VPWR VPWR DEC0.D0.AND2/X sky130_fd_sc_hd__and4bb_2
Xfill_30_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_42_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_35_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[24\].RFW.BIT\[4\].OBUF2 REGF\[24\].RFW.BIT\[4\].FF/Q REGF\[24\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[4] sky130_fd_sc_hd__ebufn_2
Xfill_39_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_39_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.BIT\[29\].OBUF1 REGF\[3\].RFW.BIT\[29\].FF/Q REGF\[3\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[29] sky130_fd_sc_hd__ebufn_2
Xfill_39_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_39_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[29\].RFW.BIT\[22\].OBUF2 REGF\[29\].RFW.BIT\[22\].FF/Q REGF\[29\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[22] sky130_fd_sc_hd__ebufn_2
Xfill_55_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_2_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_55_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_55_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_55_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_55_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_2_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_2_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[21\].RFW.BIT\[24\].OBUF1 REGF\[21\].RFW.BIT\[24\].FF/Q REGF\[21\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[24] sky130_fd_sc_hd__ebufn_2
XREGF\[6\].RFW.BIT\[14\].OBUF1 REGF\[6\].RFW.BIT\[14\].FF/Q REGF\[6\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[14] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.BIT\[20\].OBUF1 REGF\[19\].RFW.BIT\[20\].FF/Q REGF\[19\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[20] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.BIT\[0\].OBUF1 REGF\[28\].RFW.BIT\[0\].FF/Q REGF\[28\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[0] sky130_fd_sc_hd__ebufn_2
Xfill_56_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_49_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_4_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XREGF\[25\].RFW.BIT\[25\].OBUF2 REGF\[25\].RFW.BIT\[25\].FF/Q REGF\[25\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[25] sky130_fd_sc_hd__ebufn_2
XREGF\[9\].RFW.BIT\[27\].FF REGF\[9\].RFW.CG\[3\]/GCLK DW[27] VGND VGND VPWR VPWR
+ REGF\[9\].RFW.BIT\[27\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[15\].RFW.BIT\[17\].FF REGF\[15\].RFW.CG\[2\]/GCLK DW[17] VGND VGND VPWR VPWR
+ REGF\[15\].RFW.BIT\[17\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[30\].RFW.BIT\[14\].OBUF2 REGF\[30\].RFW.BIT\[14\].FF/Q REGF\[30\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[14] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[4\].OBUF2 REGF\[26\].RFW.BIT\[4\].FF/Q REGF\[26\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[4] sky130_fd_sc_hd__ebufn_2
XREGF\[2\].RFW.BIT\[17\].OBUF1 REGF\[2\].RFW.BIT\[17\].FF/Q REGF\[2\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[17] sky130_fd_sc_hd__ebufn_2
XREGF\[3\].RFW.BIT\[30\].OBUF1 REGF\[3\].RFW.BIT\[30\].FF/Q REGF\[3\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[30] sky130_fd_sc_hd__ebufn_2
Xtap_14_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[15\].RFW.BIT\[23\].OBUF1 REGF\[15\].RFW.BIT\[23\].FF/Q REGF\[15\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[23] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.BIT\[10\].OBUF2 REGF\[28\].RFW.BIT\[10\].FF/Q REGF\[28\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[10] sky130_fd_sc_hd__ebufn_2
Xtap_7_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[12\].OBUF1 REGF\[20\].RFW.BIT\[12\].FF/Q REGF\[20\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[12] sky130_fd_sc_hd__ebufn_2
Xfill_25_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_25_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_25_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_25_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_25_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_41_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_41_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_41_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDEC2.D1.ABUF\[1\] RW[1] VGND VGND VPWR VPWR DEC2.D1.AND7/B sky130_fd_sc_hd__clkbuf_2
XREGF\[26\].RFW.BIT\[27\].FF REGF\[26\].RFW.CG\[3\]/GCLK DW[27] VGND VGND VPWR VPWR
+ REGF\[26\].RFW.BIT\[27\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_41_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_41_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_41_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[21\].RFW.BIT\[28\].OBUF2 REGF\[21\].RFW.BIT\[28\].FF/Q REGF\[21\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[28] sky130_fd_sc_hd__ebufn_2
XREGF\[7\].RFW.BIT\[31\].OBUF2 REGF\[7\].RFW.BIT\[31\].FF/Q REGF\[7\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[31] sky130_fd_sc_hd__ebufn_2
XREGF\[6\].RFW.BIT\[18\].OBUF2 REGF\[6\].RFW.BIT\[18\].FF/Q REGF\[6\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[18] sky130_fd_sc_hd__ebufn_2
Xfill_42_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_35_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[19\].RFW.BIT\[24\].OBUF2 REGF\[19\].RFW.BIT\[24\].FF/Q REGF\[19\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[24] sky130_fd_sc_hd__ebufn_2
Xfill_28_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[28\].RFW.BIT\[4\].OBUF2 REGF\[28\].RFW.BIT\[4\].FF/Q REGF\[28\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[4] sky130_fd_sc_hd__ebufn_2
XREGF\[11\].RFW.BIT\[26\].OBUF1 REGF\[11\].RFW.BIT\[26\].FF/Q REGF\[11\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[26] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[13\].OBUF2 REGF\[24\].RFW.BIT\[13\].FF/Q REGF\[24\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[13] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.INV2\[1\] DEC1.D0.AND5/X VGND VGND VPWR VPWR REGF\[5\].RFW.INV2\[1\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[30\].RFW.BIT\[7\].OBUF1 REGF\[30\].RFW.BIT\[7\].FF/Q REGF\[30\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[7] sky130_fd_sc_hd__ebufn_2
XREGF\[6\].RFW.BIT\[12\].FF REGF\[6\].RFW.CG\[1\]/GCLK DW[12] VGND VGND VPWR VPWR
+ REGF\[6\].RFW.BIT\[12\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_61_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_54_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[14\].RFW.BIT\[11\].OBUF1 REGF\[14\].RFW.BIT\[11\].FF/Q REGF\[14\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[11] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.BIT\[2\].OBUF2 REGF\[21\].RFW.BIT\[2\].FF/Q REGF\[21\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[2] sky130_fd_sc_hd__ebufn_2
XREGF\[15\].RFW.BIT\[27\].OBUF2 REGF\[15\].RFW.BIT\[27\].FF/Q REGF\[15\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[27] sky130_fd_sc_hd__ebufn_2
Xfill_11_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_11_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_11_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_11_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_11_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[16\].OBUF2 REGF\[20\].RFW.BIT\[16\].FF/Q REGF\[20\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[16] sky130_fd_sc_hd__ebufn_2
XREGF\[23\].RFW.BIT\[12\].FF REGF\[23\].RFW.CG\[1\]/GCLK DW[12] VGND VGND VPWR VPWR
+ REGF\[23\].RFW.BIT\[12\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_48_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.BIT\[12\].OBUF2 REGF\[18\].RFW.BIT\[12\].FF/Q REGF\[18\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[12] sky130_fd_sc_hd__ebufn_2
Xfill_36_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_36_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[1\].RFW.INV1\[2\] DEC0.D0.AND1/X VGND VGND VPWR VPWR REGF\[1\].RFW.INV1\[2\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_36_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[10\].RFW.BIT\[14\].OBUF1 REGF\[10\].RFW.BIT\[14\].FF/Q REGF\[10\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[14] sky130_fd_sc_hd__ebufn_2
Xfill_52_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_52_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_52_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC2.D2.AND7 DEC2.D2.AND7/A DEC2.D2.AND7/B DEC2.D2.AND7/C DEC2.D2.AND7/D VGND VGND
+ VPWR VPWR DEC2.D2.AND7/X sky130_fd_sc_hd__and4_2
XREGF\[12\].RFW.BIT\[25\].FF REGF\[12\].RFW.CG\[3\]/GCLK DW[25] VGND VGND VPWR VPWR
+ REGF\[12\].RFW.BIT\[25\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_8_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfill_8_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_8_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[23\].RFW.BIT\[2\].OBUF2 REGF\[23\].RFW.BIT\[2\].FF/Q REGF\[23\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[2] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.INV1\[0\] DEC0.D2.AND5/X VGND VGND VPWR VPWR REGF\[21\].RFW.INV1\[0\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_40_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_33_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_26_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_19_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[2\].RFW.BIT\[22\].OBUF2 REGF\[2\].RFW.BIT\[22\].FF/Q REGF\[2\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[22] sky130_fd_sc_hd__ebufn_2
XREGF\[6\].RFW.CGAND DEC2.D0.AND6/X WE VGND VGND VPWR VPWR REGF\[6\].RFW.CGAND/X sky130_fd_sc_hd__and2_1
XREGF\[14\].RFW.BIT\[15\].OBUF2 REGF\[14\].RFW.BIT\[15\].FF/Q REGF\[14\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[15] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.CG\[3\] CLK REGF\[28\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[28\].RFW.CG\[3\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_22_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_22_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_22_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[25\].RFW.BIT\[2\].OBUF2 REGF\[25\].RFW.BIT\[2\].FF/Q REGF\[25\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[2] sky130_fd_sc_hd__ebufn_2
XREGF\[7\].RFW.BIT\[18\].FF REGF\[7\].RFW.CG\[2\]/GCLK DW[18] VGND VGND VPWR VPWR
+ REGF\[7\].RFW.BIT\[18\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[11\].RFW.BIT\[31\].OBUF2 REGF\[11\].RFW.BIT\[31\].FF/Q REGF\[11\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[31] sky130_fd_sc_hd__ebufn_2
XREGF\[10\].RFW.BIT\[18\].OBUF2 REGF\[10\].RFW.BIT\[18\].FF/Q REGF\[10\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[18] sky130_fd_sc_hd__ebufn_2
XREGF\[3\].RFW.BIT\[20\].FF REGF\[3\].RFW.CG\[2\]/GCLK DW[20] VGND VGND VPWR VPWR
+ REGF\[3\].RFW.BIT\[20\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[1\].RFW.CG\[1\] CLK REGF\[1\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[1\].RFW.CG\[1\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XDEC1.D2.ABUF\[2\] RB[2] VGND VGND VPWR VPWR DEC1.D2.AND7/C sky130_fd_sc_hd__clkbuf_2
Xfill_47_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_47_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_47_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_47_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_47_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_47_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[1\].RFW.BIT\[10\].OBUF2 REGF\[1\].RFW.BIT\[10\].FF/Q REGF\[1\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[10] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[28\].OBUF1 REGF\[26\].RFW.BIT\[28\].FF/Q REGF\[26\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[28] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.CG\[0\] CLK REGF\[27\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[27\].RFW.CG\[0\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[31\].RFW.BIT\[17\].OBUF1 REGF\[31\].RFW.BIT\[17\].FF/Q REGF\[31\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[17] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.INV1\[1\] DEC0.D2.AND0/Y VGND VGND VPWR VPWR REGF\[16\].RFW.INV1\[1\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[24\].RFW.BIT\[18\].FF REGF\[24\].RFW.CG\[2\]/GCLK DW[18] VGND VGND VPWR VPWR
+ REGF\[24\].RFW.BIT\[18\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[20\].RFW.BIT\[20\].FF REGF\[20\].RFW.CG\[2\]/GCLK DW[20] VGND VGND VPWR VPWR
+ REGF\[20\].RFW.BIT\[20\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[29\].RFW.BIT\[13\].OBUF1 REGF\[29\].RFW.BIT\[13\].FF/Q REGF\[29\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[13] sky130_fd_sc_hd__ebufn_2
Xfill_31_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XREGF\[27\].RFW.BIT\[2\].OBUF2 REGF\[27\].RFW.BIT\[2\].FF/Q REGF\[27\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[2] sky130_fd_sc_hd__ebufn_2
Xfill_24_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_17_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.INV2\[2\] DEC1.D3.AND7/X VGND VGND VPWR VPWR REGF\[31\].RFW.INV2\[2\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[19\].RFW.BIT\[25\].FF REGF\[19\].RFW.CG\[3\]/GCLK DW[25] VGND VGND VPWR VPWR
+ REGF\[19\].RFW.BIT\[25\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_46_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.BIT\[30\].FF REGF\[31\].RFW.CG\[3\]/GCLK DW[30] VGND VGND VPWR VPWR
+ REGF\[31\].RFW.BIT\[30\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[16\].RFW.CG\[3\] CLK REGF\[16\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[16\].RFW.CG\[3\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[20\].RFW.BIT\[0\].OBUF2 REGF\[20\].RFW.BIT\[0\].FF/Q REGF\[20\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[0] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.CGAND DEC2.D2.AND0/Y WE VGND VGND VPWR VPWR REGF\[16\].RFW.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_17_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_17_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_17_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_17_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_17_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_33_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[25\].RFW.BIT\[16\].OBUF1 REGF\[25\].RFW.BIT\[16\].FF/Q REGF\[25\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[16] sky130_fd_sc_hd__ebufn_2
Xfill_33_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDEC0.D3.AND0 DEC0.D3.AND7/A DEC0.D3.AND7/B DEC0.D3.AND7/C DEC0.D3.AND7/D VGND VGND
+ VPWR VPWR DEC0.D3.AND0/Y sky130_fd_sc_hd__nor4b_2
XREGF\[29\].RFW.BIT\[2\].OBUF2 REGF\[29\].RFW.BIT\[2\].FF/Q REGF\[29\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[2] sky130_fd_sc_hd__ebufn_2
Xfill_58_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_58_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_5_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_5_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_5_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_5_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_5_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_10_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_8_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[15\].RFW.CG\[0\] CLK REGF\[15\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[15\].RFW.CG\[0\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[31\].RFW.BIT\[5\].OBUF1 REGF\[31\].RFW.BIT\[5\].FF/Q REGF\[31\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[5] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.BIT\[17\].OBUF2 REGF\[29\].RFW.BIT\[17\].FF/Q REGF\[29\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[17] sky130_fd_sc_hd__ebufn_2
XREGF\[10\].RFW.BIT\[16\].FF REGF\[10\].RFW.CG\[2\]/GCLK DW[16] VGND VGND VPWR VPWR
+ REGF\[10\].RFW.BIT\[16\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[21\].RFW.BIT\[19\].OBUF1 REGF\[21\].RFW.BIT\[19\].FF/Q REGF\[21\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[19] sky130_fd_sc_hd__ebufn_2
XREGF\[22\].RFW.BIT\[0\].OBUF2 REGF\[22\].RFW.BIT\[0\].FF/Q REGF\[22\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[0] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.BIT\[26\].FF REGF\[4\].RFW.CG\[3\]/GCLK DW[26] VGND VGND VPWR VPWR
+ REGF\[4\].RFW.BIT\[26\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[10\].RFW.INV2\[2\] DEC1.D1.AND2/X VGND VGND VPWR VPWR REGF\[10\].RFW.INV2\[2\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[16\].RFW.BIT\[10\].FF REGF\[16\].RFW.CG\[1\]/GCLK DW[10] VGND VGND VPWR VPWR
+ REGF\[16\].RFW.BIT\[10\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[7\].RFW.BIT\[22\].OBUF1 REGF\[7\].RFW.BIT\[22\].FF/Q REGF\[7\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[22] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.INV2\[3\] DEC1.D3.AND2/X VGND VGND VPWR VPWR REGF\[26\].RFW.INV2\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[19\].RFW.BIT\[15\].OBUF1 REGF\[19\].RFW.BIT\[15\].FF/Q REGF\[19\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[15] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.BIT\[9\].FF REGF\[19\].RFW.CG\[1\]/GCLK DW[9] VGND VGND VPWR VPWR
+ REGF\[19\].RFW.BIT\[9\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_44_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[21\].RFW.BIT\[26\].FF REGF\[21\].RFW.CG\[3\]/GCLK DW[26] VGND VGND VPWR VPWR
+ REGF\[21\].RFW.BIT\[26\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_56_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_28_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_28_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[27\].RFW.BIT\[20\].FF REGF\[27\].RFW.CG\[2\]/GCLK DW[20] VGND VGND VPWR VPWR
+ REGF\[27\].RFW.BIT\[20\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_28_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.BIT\[22\].OBUF2 REGF\[31\].RFW.BIT\[22\].FF/Q REGF\[31\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[22] sky130_fd_sc_hd__ebufn_2
Xfill_44_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_44_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_44_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.BIT\[25\].OBUF1 REGF\[3\].RFW.BIT\[25\].FF/Q REGF\[3\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[25] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[0\].OBUF2 REGF\[24\].RFW.BIT\[0\].FF/Q REGF\[24\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[0] sky130_fd_sc_hd__ebufn_2
Xfill_60_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_60_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_60_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[15\].RFW.BIT\[18\].OBUF1 REGF\[15\].RFW.BIT\[18\].FF/Q REGF\[15\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[18] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[31\].OBUF1 REGF\[16\].RFW.BIT\[31\].FF/Q REGF\[16\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[31] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.BIT\[20\].OBUF1 REGF\[21\].RFW.BIT\[20\].FF/Q REGF\[21\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[20] sky130_fd_sc_hd__ebufn_2
XREGF\[31\].RFW.BIT\[9\].OBUF2 REGF\[31\].RFW.BIT\[9\].FF/Q REGF\[31\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[9] sky130_fd_sc_hd__ebufn_2
Xfill_58_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[1\].RFW.BIT\[11\].FF REGF\[1\].RFW.CG\[1\]/GCLK DW[11] VGND VGND VPWR VPWR
+ REGF\[1\].RFW.BIT\[11\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xgenblk1.RFW0.INV1\[2\] DEC0.D0.AND0/Y VGND VGND VPWR VPWR genblk1.RFW0.INV1\[2\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[6\].RFW.BIT\[10\].OBUF1 REGF\[6\].RFW.BIT\[10\].FF/Q REGF\[6\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[10] sky130_fd_sc_hd__ebufn_2
Xfill_6_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[7\].RFW.BIT\[26\].OBUF2 REGF\[7\].RFW.BIT\[26\].FF/Q REGF\[7\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[26] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.BIT\[19\].OBUF2 REGF\[19\].RFW.BIT\[19\].FF/Q REGF\[19\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[19] sky130_fd_sc_hd__ebufn_2
Xtap_16_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[25\].RFW.BIT\[21\].OBUF2 REGF\[25\].RFW.BIT\[21\].FF/Q REGF\[25\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[21] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[0\].OBUF2 REGF\[26\].RFW.BIT\[0\].FF/Q REGF\[26\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[0] sky130_fd_sc_hd__ebufn_2
XREGF\[30\].RFW.BIT\[10\].OBUF2 REGF\[30\].RFW.BIT\[10\].FF/Q REGF\[30\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[10] sky130_fd_sc_hd__ebufn_2
XREGF\[2\].RFW.BIT\[13\].OBUF1 REGF\[2\].RFW.BIT\[13\].FF/Q REGF\[2\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[13] sky130_fd_sc_hd__ebufn_2
Xfill_14_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_14_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_14_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_30_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_30_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDEC0.D0.AND3 DEC0.D0.AND7/C DEC0.D0.AND7/B DEC0.D0.AND7/A DEC0.D0.AND7/D VGND VGND
+ VPWR VPWR DEC0.D0.AND3/X sky130_fd_sc_hd__and4b_2
Xfill_30_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_42_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_35_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[17\].RFW.BIT\[16\].FF REGF\[17\].RFW.CG\[2\]/GCLK DW[16] VGND VGND VPWR VPWR
+ REGF\[17\].RFW.BIT\[16\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_39_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_39_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[3\].RFW.BIT\[29\].OBUF2 REGF\[3\].RFW.BIT\[29\].FF/Q REGF\[3\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[29] sky130_fd_sc_hd__ebufn_2
Xfill_39_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_39_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_55_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_55_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_55_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_55_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_55_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_2_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_2_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_55_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[21\].RFW.BIT\[24\].OBUF2 REGF\[21\].RFW.BIT\[24\].FF/Q REGF\[21\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[24] sky130_fd_sc_hd__ebufn_2
XREGF\[6\].RFW.BIT\[14\].OBUF2 REGF\[6\].RFW.BIT\[14\].FF/Q REGF\[6\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[14] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.BIT\[20\].OBUF2 REGF\[19\].RFW.BIT\[20\].FF/Q REGF\[19\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[20] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.BIT\[0\].OBUF2 REGF\[28\].RFW.BIT\[0\].FF/Q REGF\[28\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[0] sky130_fd_sc_hd__ebufn_2
XREGF\[11\].RFW.BIT\[22\].OBUF1 REGF\[11\].RFW.BIT\[22\].FF/Q REGF\[11\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[22] sky130_fd_sc_hd__ebufn_2
Xfill_56_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[28\].RFW.BIT\[26\].FF REGF\[28\].RFW.CG\[3\]/GCLK DW[26] VGND VGND VPWR VPWR
+ REGF\[28\].RFW.BIT\[26\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_49_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[30\].RFW.BIT\[3\].OBUF1 REGF\[30\].RFW.BIT\[3\].FF/Q REGF\[30\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[3] sky130_fd_sc_hd__ebufn_2
Xfill_4_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[2\].RFW.BIT\[17\].FF REGF\[2\].RFW.CG\[2\]/GCLK DW[17] VGND VGND VPWR VPWR
+ REGF\[2\].RFW.BIT\[17\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[2\].RFW.BIT\[17\].OBUF2 REGF\[2\].RFW.BIT\[17\].FF/Q REGF\[2\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[17] sky130_fd_sc_hd__ebufn_2
XREGF\[3\].RFW.BIT\[30\].OBUF2 REGF\[3\].RFW.BIT\[30\].FF/Q REGF\[3\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[30] sky130_fd_sc_hd__ebufn_2
Xtap_14_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[15\].RFW.BIT\[23\].OBUF2 REGF\[15\].RFW.BIT\[23\].FF/Q REGF\[15\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[23] sky130_fd_sc_hd__ebufn_2
XREGF\[8\].RFW.BIT\[11\].FF REGF\[8\].RFW.CG\[1\]/GCLK DW[11] VGND VGND VPWR VPWR
+ REGF\[8\].RFW.BIT\[11\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_7_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[12\].OBUF2 REGF\[20\].RFW.BIT\[12\].FF/Q REGF\[20\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[12] sky130_fd_sc_hd__ebufn_2
Xfill_25_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_25_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_25_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_25_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_41_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_41_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_41_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_41_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_41_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[10\].RFW.BIT\[10\].OBUF1 REGF\[10\].RFW.BIT\[10\].FF/Q REGF\[10\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[10] sky130_fd_sc_hd__ebufn_2
XREGF\[8\].RFW.INV2\[2\] DEC1.D1.AND0/Y VGND VGND VPWR VPWR REGF\[8\].RFW.INV2\[2\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_35_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[25\].RFW.BIT\[11\].FF REGF\[25\].RFW.CG\[1\]/GCLK DW[11] VGND VGND VPWR VPWR
+ REGF\[25\].RFW.BIT\[11\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_28_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[11\].RFW.BIT\[26\].OBUF2 REGF\[11\].RFW.BIT\[26\].FF/Q REGF\[11\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[26] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.CGAND DEC2.D0.AND5/X WE VGND VGND VPWR VPWR REGF\[5\].RFW.CGAND/X sky130_fd_sc_hd__and2_1
XREGF\[28\].RFW.INV2\[0\] DEC1.D3.AND4/X VGND VGND VPWR VPWR REGF\[28\].RFW.INV2\[0\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[30\].RFW.BIT\[7\].OBUF2 REGF\[30\].RFW.BIT\[7\].FF/Q REGF\[30\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[7] sky130_fd_sc_hd__ebufn_2
Xfill_61_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_54_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[14\].RFW.BIT\[11\].OBUF2 REGF\[14\].RFW.BIT\[11\].FF/Q REGF\[14\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[11] sky130_fd_sc_hd__ebufn_2
XREGF\[14\].RFW.BIT\[24\].FF REGF\[14\].RFW.CG\[3\]/GCLK DW[24] VGND VGND VPWR VPWR
+ REGF\[14\].RFW.BIT\[24\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[30\].RFW.BIT\[27\].FF REGF\[30\].RFW.CG\[3\]/GCLK DW[27] VGND VGND VPWR VPWR
+ REGF\[30\].RFW.BIT\[27\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_47_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_2_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[24\].RFW.CG\[2\] CLK REGF\[24\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[24\].RFW.CG\[2\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[17\].RFW.BIT\[0\].FF REGF\[17\].RFW.CG\[0\]/GCLK DW[0] VGND VGND VPWR VPWR
+ REGF\[17\].RFW.BIT\[0\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[4\].RFW.INV1\[3\] DEC0.D0.AND4/X VGND VGND VPWR VPWR REGF\[4\].RFW.INV1\[3\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_11_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_11_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_11_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_11_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_11_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xtap_12_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_5_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_36_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[16\].RFW.BIT\[2\].FF REGF\[16\].RFW.CG\[0\]/GCLK DW[2] VGND VGND VPWR VPWR
+ REGF\[16\].RFW.BIT\[2\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_36_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_36_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[10\].RFW.BIT\[14\].OBUF2 REGF\[10\].RFW.BIT\[14\].FF/Q REGF\[10\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[14] sky130_fd_sc_hd__ebufn_2
Xfill_52_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_52_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_52_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[24\].RFW.INV1\[1\] DEC0.D3.AND0/Y VGND VGND VPWR VPWR REGF\[24\].RFW.INV1\[1\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[8\].RFW.BIT\[29\].OBUF1 REGF\[8\].RFW.BIT\[29\].FF/Q REGF\[8\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[29] sky130_fd_sc_hd__ebufn_2
Xfill_8_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_8_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[15\].RFW.BIT\[4\].FF REGF\[15\].RFW.CG\[0\]/GCLK DW[4] VGND VGND VPWR VPWR
+ REGF\[15\].RFW.BIT\[4\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[26\].RFW.BIT\[24\].OBUF1 REGF\[26\].RFW.BIT\[24\].FF/Q REGF\[26\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[24] sky130_fd_sc_hd__ebufn_2
XREGF\[9\].RFW.BIT\[17\].FF REGF\[9\].RFW.CG\[2\]/GCLK DW[17] VGND VGND VPWR VPWR
+ REGF\[9\].RFW.BIT\[17\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_40_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_33_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.BIT\[13\].OBUF1 REGF\[31\].RFW.BIT\[13\].FF/Q REGF\[31\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[13] sky130_fd_sc_hd__ebufn_2
Xfill_26_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_19_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[14\].RFW.BIT\[6\].FF REGF\[14\].RFW.CG\[0\]/GCLK DW[6] VGND VGND VPWR VPWR
+ REGF\[14\].RFW.BIT\[6\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[12\].RFW.CG\[2\] CLK REGF\[12\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[12\].RFW.CG\[2\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[15\].RFW.CGAND DEC2.D1.AND7/X WE VGND VGND VPWR VPWR REGF\[15\].RFW.CGAND/X
+ sky130_fd_sc_hd__and2_1
XREGF\[26\].RFW.BIT\[17\].FF REGF\[26\].RFW.CG\[2\]/GCLK DW[17] VGND VGND VPWR VPWR
+ REGF\[26\].RFW.BIT\[17\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[29\].RFW.BIT\[2\].FF REGF\[29\].RFW.CG\[0\]/GCLK DW[2] VGND VGND VPWR VPWR
+ REGF\[29\].RFW.BIT\[2\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[13\].RFW.BIT\[8\].FF REGF\[13\].RFW.CG\[1\]/GCLK DW[8] VGND VGND VPWR VPWR
+ REGF\[13\].RFW.BIT\[8\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[22\].RFW.BIT\[27\].OBUF1 REGF\[22\].RFW.BIT\[27\].FF/Q REGF\[22\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[27] sky130_fd_sc_hd__ebufn_2
Xfill_22_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_22_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[7\].RFW.BIT\[17\].OBUF1 REGF\[7\].RFW.BIT\[17\].FF/Q REGF\[7\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[17] sky130_fd_sc_hd__ebufn_2
Xfill_22_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[8\].RFW.BIT\[30\].OBUF1 REGF\[8\].RFW.BIT\[30\].FF/Q REGF\[8\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[30] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.BIT\[4\].FF REGF\[28\].RFW.CG\[0\]/GCLK DW[4] VGND VGND VPWR VPWR
+ REGF\[28\].RFW.BIT\[4\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_10_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[25\].RFW.BIT\[12\].OBUF1 REGF\[25\].RFW.BIT\[12\].FF/Q REGF\[25\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[12] sky130_fd_sc_hd__ebufn_2
Xfill_47_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_47_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_47_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_47_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_47_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_47_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[19\].RFW.INV1\[2\] DEC0.D2.AND3/X VGND VGND VPWR VPWR REGF\[19\].RFW.INV1\[2\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[27\].RFW.BIT\[6\].FF REGF\[27\].RFW.CG\[0\]/GCLK DW[6] VGND VGND VPWR VPWR
+ REGF\[27\].RFW.BIT\[6\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[26\].RFW.BIT\[28\].OBUF2 REGF\[26\].RFW.BIT\[28\].FF/Q REGF\[26\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[28] sky130_fd_sc_hd__ebufn_2
XREGF\[31\].RFW.BIT\[17\].OBUF2 REGF\[31\].RFW.BIT\[17\].FF/Q REGF\[31\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[17] sky130_fd_sc_hd__ebufn_2
XREGF\[31\].RFW.BIT\[1\].OBUF1 REGF\[31\].RFW.BIT\[1\].FF/Q REGF\[31\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[1] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[26\].OBUF1 REGF\[16\].RFW.BIT\[26\].FF/Q REGF\[16\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[26] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.BIT\[13\].OBUF2 REGF\[29\].RFW.BIT\[13\].FF/Q REGF\[29\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[13] sky130_fd_sc_hd__ebufn_2
Xfill_31_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[26\].RFW.BIT\[8\].FF REGF\[26\].RFW.CG\[1\]/GCLK DW[8] VGND VGND VPWR VPWR
+ REGF\[26\].RFW.BIT\[8\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_24_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_17_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[21\].RFW.BIT\[15\].OBUF1 REGF\[21\].RFW.BIT\[15\].FF/Q REGF\[21\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[15] sky130_fd_sc_hd__ebufn_2
XDEC1.D0.ABUF\[1\] RB[1] VGND VGND VPWR VPWR DEC1.D0.AND7/B sky130_fd_sc_hd__clkbuf_2
XREGF\[19\].RFW.BIT\[11\].OBUF1 REGF\[19\].RFW.BIT\[11\].FF/Q REGF\[19\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[11] sky130_fd_sc_hd__ebufn_2
Xtap_46_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.BIT\[25\].FF REGF\[6\].RFW.CG\[3\]/GCLK DW[25] VGND VGND VPWR VPWR
+ REGF\[6\].RFW.BIT\[25\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[12\].RFW.BIT\[15\].FF REGF\[12\].RFW.CG\[1\]/GCLK DW[15] VGND VGND VPWR VPWR
+ REGF\[12\].RFW.BIT\[15\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_17_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_17_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_17_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_17_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_17_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.BIT\[29\].OBUF1 REGF\[12\].RFW.BIT\[29\].FF/Q REGF\[12\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[29] sky130_fd_sc_hd__ebufn_2
Xfill_33_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_33_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[25\].RFW.BIT\[16\].OBUF2 REGF\[25\].RFW.BIT\[16\].FF/Q REGF\[25\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[16] sky130_fd_sc_hd__ebufn_2
Xfill_33_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_33_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_58_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC0.D3.AND1 DEC0.D3.AND7/C DEC0.D3.AND7/B DEC0.D3.AND7/A DEC0.D3.AND7/D VGND VGND
+ VPWR VPWR DEC0.D3.AND1/X sky130_fd_sc_hd__and4bb_2
Xfill_58_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_58_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_58_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_5_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.BIT\[21\].OBUF1 REGF\[3\].RFW.BIT\[21\].FF/Q REGF\[3\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[21] sky130_fd_sc_hd__ebufn_2
Xfill_5_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_5_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_5_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[15\].RFW.BIT\[14\].OBUF1 REGF\[15\].RFW.BIT\[14\].FF/Q REGF\[15\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[14] sky130_fd_sc_hd__ebufn_2
XREGF\[23\].RFW.BIT\[25\].FF REGF\[23\].RFW.CG\[3\]/GCLK DW[25] VGND VGND VPWR VPWR
+ REGF\[23\].RFW.BIT\[25\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_10_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[13\].RFW.INV2\[3\] DEC1.D1.AND5/X VGND VGND VPWR VPWR REGF\[13\].RFW.INV2\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[31\].RFW.BIT\[5\].OBUF2 REGF\[31\].RFW.BIT\[5\].FF/Q REGF\[31\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[5] sky130_fd_sc_hd__ebufn_2
XREGF\[9\].RFW.BIT\[9\].FF REGF\[9\].RFW.CG\[1\]/GCLK DW[9] VGND VGND VPWR VPWR REGF\[9\].RFW.BIT\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[21\].RFW.BIT\[19\].OBUF2 REGF\[21\].RFW.BIT\[19\].FF/Q REGF\[21\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[19] sky130_fd_sc_hd__ebufn_2
XREGF\[7\].RFW.BIT\[22\].OBUF2 REGF\[7\].RFW.BIT\[22\].FF/Q REGF\[7\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[22] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.BIT\[15\].OBUF2 REGF\[19\].RFW.BIT\[15\].FF/Q REGF\[19\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[15] sky130_fd_sc_hd__ebufn_2
XREGF\[6\].RFW.INV1\[0\] DEC0.D0.AND6/X VGND VGND VPWR VPWR REGF\[6\].RFW.INV1\[0\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[3\].RFW.BIT\[10\].FF REGF\[3\].RFW.CG\[1\]/GCLK DW[10] VGND VGND VPWR VPWR
+ REGF\[3\].RFW.BIT\[10\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[12\].RFW.BIT\[30\].OBUF1 REGF\[12\].RFW.BIT\[30\].FF/Q REGF\[12\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[30] sky130_fd_sc_hd__ebufn_2
XREGF\[11\].RFW.BIT\[17\].OBUF1 REGF\[11\].RFW.BIT\[17\].FF/Q REGF\[11\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[17] sky130_fd_sc_hd__ebufn_2
Xtap_44_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_28_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_28_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_28_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_44_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_44_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_44_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgenblk1.RFW0.BIT\[31\].OBUF1 genblk1.RFW0.TIE\[3\]/LO genblk1.RFW0.INV1\[3\]/Y VGND
+ VGND VPWR VPWR DA[31] sky130_fd_sc_hd__ebufn_2
XREGF\[20\].RFW.BIT\[10\].FF REGF\[20\].RFW.CG\[1\]/GCLK DW[10] VGND VGND VPWR VPWR
+ REGF\[20\].RFW.BIT\[10\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[3\].RFW.BIT\[25\].OBUF2 REGF\[3\].RFW.BIT\[25\].FF/Q REGF\[3\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[25] sky130_fd_sc_hd__ebufn_2
Xfill_60_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_60_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[15\].RFW.BIT\[18\].OBUF2 REGF\[15\].RFW.BIT\[18\].FF/Q REGF\[15\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[18] sky130_fd_sc_hd__ebufn_2
Xfill_60_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[16\].RFW.BIT\[31\].OBUF2 REGF\[16\].RFW.BIT\[31\].FF/Q REGF\[16\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[31] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.BIT\[20\].OBUF2 REGF\[21\].RFW.BIT\[20\].FF/Q REGF\[21\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[20] sky130_fd_sc_hd__ebufn_2
Xfill_58_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.BIT\[10\].OBUF2 REGF\[6\].RFW.BIT\[10\].FF/Q REGF\[6\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[10] sky130_fd_sc_hd__ebufn_2
Xfill_6_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[19\].RFW.BIT\[15\].FF REGF\[19\].RFW.CG\[1\]/GCLK DW[15] VGND VGND VPWR VPWR
+ REGF\[19\].RFW.BIT\[15\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[31\].RFW.BIT\[20\].FF REGF\[31\].RFW.CG\[2\]/GCLK DW[20] VGND VGND VPWR VPWR
+ REGF\[31\].RFW.BIT\[20\].FF/Q sky130_fd_sc_hd__dfxtp_1
XDEC0.D1.ABUF\[2\] RA[2] VGND VGND VPWR VPWR DEC0.D1.AND7/C sky130_fd_sc_hd__clkbuf_2
XREGF\[2\].RFW.BIT\[13\].OBUF2 REGF\[2\].RFW.BIT\[13\].FF/Q REGF\[2\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[13] sky130_fd_sc_hd__ebufn_2
Xfill_14_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_14_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_30_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XDEC0.D0.AND4 DEC0.D0.AND7/A DEC0.D0.AND7/B DEC0.D0.AND7/C DEC0.D0.AND7/D VGND VGND
+ VPWR VPWR DEC0.D0.AND4/X sky130_fd_sc_hd__and4bb_2
Xfill_30_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_30_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_42_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_35_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[10\].RFW.BIT\[1\].FF REGF\[10\].RFW.CG\[0\]/GCLK DW[1] VGND VGND VPWR VPWR
+ REGF\[10\].RFW.BIT\[1\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_28_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_39_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_55_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_55_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_55_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_55_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_55_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_2_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_2_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_55_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[4\].RFW.BIT\[16\].FF REGF\[4\].RFW.CG\[2\]/GCLK DW[16] VGND VGND VPWR VPWR
+ REGF\[4\].RFW.BIT\[16\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[4\].RFW.CGAND DEC2.D0.AND4/X WE VGND VGND VPWR VPWR REGF\[4\].RFW.CGAND/X sky130_fd_sc_hd__and2_1
XDEC1.TIE VGND VGND VPWR VPWR DEC1.TIE/HI DEC1.TIE/LO sky130_fd_sc_hd__conb_1
XREGF\[11\].RFW.BIT\[22\].OBUF2 REGF\[11\].RFW.BIT\[22\].FF/Q REGF\[11\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[22] sky130_fd_sc_hd__ebufn_2
Xfill_56_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_49_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[9\].RFW.CG\[1\] CLK REGF\[9\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[9\].RFW.CG\[1\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[20\].RFW.CG\[1\] CLK REGF\[20\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[20\].RFW.CG\[1\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[30\].RFW.BIT\[3\].OBUF2 REGF\[30\].RFW.BIT\[3\].FF/Q REGF\[30\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[3] sky130_fd_sc_hd__ebufn_2
Xfill_4_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[21\].RFW.BIT\[16\].FF REGF\[21\].RFW.CG\[2\]/GCLK DW[16] VGND VGND VPWR VPWR
+ REGF\[21\].RFW.BIT\[16\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[26\].RFW.BIT\[19\].OBUF1 REGF\[26\].RFW.BIT\[19\].FF/Q REGF\[26\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[19] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[10\].FF REGF\[27\].RFW.CG\[1\]/GCLK DW[10] VGND VGND VPWR VPWR
+ REGF\[27\].RFW.BIT\[10\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[23\].RFW.BIT\[1\].FF REGF\[23\].RFW.CG\[0\]/GCLK DW[1] VGND VGND VPWR VPWR
+ REGF\[23\].RFW.BIT\[1\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_14_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[10\].RFW.BIT\[29\].FF REGF\[10\].RFW.CG\[3\]/GCLK DW[29] VGND VGND VPWR VPWR
+ REGF\[10\].RFW.BIT\[29\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[16\].RFW.BIT\[23\].FF REGF\[16\].RFW.CG\[2\]/GCLK DW[23] VGND VGND VPWR VPWR
+ REGF\[16\].RFW.BIT\[23\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_25_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_25_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_25_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_25_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_25_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[22\].RFW.BIT\[3\].FF REGF\[22\].RFW.CG\[0\]/GCLK DW[3] VGND VGND VPWR VPWR
+ REGF\[22\].RFW.BIT\[3\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_41_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_41_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_41_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_41_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_41_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC1.D.AND0 RB[3] RB[4] DEC1.TIE/HI VGND VGND VPWR VPWR DEC1.D.AND0/Y sky130_fd_sc_hd__nor3b_4
Xtap_40_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[10\].RFW.BIT\[10\].OBUF2 REGF\[10\].RFW.BIT\[10\].FF/Q REGF\[10\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[10] sky130_fd_sc_hd__ebufn_2
XREGF\[15\].RFW.INV2\[0\] DEC1.D1.AND7/X VGND VGND VPWR VPWR REGF\[15\].RFW.INV2\[0\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[21\].RFW.BIT\[5\].FF REGF\[21\].RFW.CG\[0\]/GCLK DW[5] VGND VGND VPWR VPWR
+ REGF\[21\].RFW.BIT\[5\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[8\].RFW.BIT\[25\].OBUF1 REGF\[8\].RFW.BIT\[25\].FF/Q REGF\[8\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[25] sky130_fd_sc_hd__ebufn_2
Xfill_28_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[26\].RFW.BIT\[20\].OBUF1 REGF\[26\].RFW.BIT\[20\].FF/Q REGF\[26\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[20] sky130_fd_sc_hd__ebufn_2
XREGF\[7\].RFW.BIT\[0\].FF REGF\[7\].RFW.CG\[0\]/GCLK DW[0] VGND VGND VPWR VPWR REGF\[7\].RFW.BIT\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[20\].RFW.BIT\[7\].FF REGF\[20\].RFW.CG\[0\]/GCLK DW[7] VGND VGND VPWR VPWR
+ REGF\[20\].RFW.BIT\[7\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_61_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_54_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[14\].RFW.CGAND DEC2.D1.AND6/X WE VGND VGND VPWR VPWR REGF\[14\].RFW.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_47_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_3_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC2.D3.ABUF\[0\] RW[0] VGND VGND VPWR VPWR DEC2.D3.AND7/A sky130_fd_sc_hd__clkbuf_2
XREGF\[6\].RFW.BIT\[2\].FF REGF\[6\].RFW.CG\[0\]/GCLK DW[2] VGND VGND VPWR VPWR REGF\[6\].RFW.BIT\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xfill_2_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[1\].RFW.BIT\[24\].FF REGF\[1\].RFW.CG\[3\]/GCLK DW[24] VGND VGND VPWR VPWR
+ REGF\[1\].RFW.BIT\[24\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[4\].RFW.BIT\[28\].OBUF1 REGF\[4\].RFW.BIT\[28\].FF/Q REGF\[4\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[28] sky130_fd_sc_hd__ebufn_2
Xfill_11_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[11\].RFW.INV1\[1\] DEC0.D1.AND3/X VGND VGND VPWR VPWR REGF\[11\].RFW.INV1\[1\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_11_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_11_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_11_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[22\].RFW.BIT\[23\].OBUF1 REGF\[22\].RFW.BIT\[23\].FF/Q REGF\[22\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[23] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.INV1\[2\] DEC0.D3.AND3/X VGND VGND VPWR VPWR REGF\[27\].RFW.INV1\[2\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[5\].RFW.BIT\[4\].FF REGF\[5\].RFW.CG\[0\]/GCLK DW[4] VGND VGND VPWR VPWR REGF\[5\].RFW.BIT\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xtap_12_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[7\].RFW.BIT\[13\].OBUF1 REGF\[7\].RFW.BIT\[13\].FF/Q REGF\[7\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[13] sky130_fd_sc_hd__ebufn_2
Xtap_5_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_36_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_36_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_36_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_52_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_52_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_52_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[28\].RFW.BIT\[16\].FF REGF\[28\].RFW.CG\[2\]/GCLK DW[16] VGND VGND VPWR VPWR
+ REGF\[28\].RFW.BIT\[16\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[8\].RFW.BIT\[29\].OBUF2 REGF\[8\].RFW.BIT\[29\].FF/Q REGF\[8\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[29] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.BIT\[6\].FF REGF\[4\].RFW.CG\[0\]/GCLK DW[6] VGND VGND VPWR VPWR REGF\[4\].RFW.BIT\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xfill_8_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_8_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[26\].RFW.BIT\[24\].OBUF2 REGF\[26\].RFW.BIT\[24\].FF/Q REGF\[26\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[24] sky130_fd_sc_hd__ebufn_2
Xfill_40_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_26_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[31\].RFW.BIT\[13\].OBUF2 REGF\[31\].RFW.BIT\[13\].FF/Q REGF\[31\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[13] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.BIT\[29\].FF REGF\[17\].RFW.CG\[3\]/GCLK DW[29] VGND VGND VPWR VPWR
+ REGF\[17\].RFW.BIT\[29\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_19_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[13\].RFW.BIT\[31\].FF REGF\[13\].RFW.CG\[3\]/GCLK DW[31] VGND VGND VPWR VPWR
+ REGF\[13\].RFW.BIT\[31\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[3\].RFW.BIT\[8\].FF REGF\[3\].RFW.CG\[1\]/GCLK DW[8] VGND VGND VPWR VPWR REGF\[3\].RFW.BIT\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[3\].RFW.BIT\[16\].OBUF1 REGF\[3\].RFW.BIT\[16\].FF/Q REGF\[3\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[16] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[22\].OBUF1 REGF\[16\].RFW.BIT\[22\].FF/Q REGF\[16\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[22] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.BIT\[11\].OBUF1 REGF\[21\].RFW.BIT\[11\].FF/Q REGF\[21\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[11] sky130_fd_sc_hd__ebufn_2
XREGF\[22\].RFW.BIT\[27\].OBUF2 REGF\[22\].RFW.BIT\[27\].FF/Q REGF\[22\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[27] sky130_fd_sc_hd__ebufn_2
Xfill_22_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_22_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[7\].RFW.BIT\[17\].OBUF2 REGF\[7\].RFW.BIT\[17\].FF/Q REGF\[7\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[17] sky130_fd_sc_hd__ebufn_2
Xfill_22_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[8\].RFW.BIT\[30\].OBUF2 REGF\[8\].RFW.BIT\[30\].FF/Q REGF\[8\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[30] sky130_fd_sc_hd__ebufn_2
Xtap_10_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.BIT\[25\].OBUF1 REGF\[12\].RFW.BIT\[25\].FF/Q REGF\[12\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[25] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.INV2\[3\] DEC1.D2.AND5/X VGND VGND VPWR VPWR REGF\[21\].RFW.INV2\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[25\].RFW.BIT\[12\].OBUF2 REGF\[25\].RFW.BIT\[12\].FF/Q REGF\[25\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[12] sky130_fd_sc_hd__ebufn_2
Xfill_47_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_47_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_47_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_47_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_47_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xtap_3_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[8\].RFW.BIT\[24\].FF REGF\[8\].RFW.CG\[3\]/GCLK DW[24] VGND VGND VPWR VPWR
+ REGF\[8\].RFW.BIT\[24\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[14\].RFW.BIT\[14\].FF REGF\[14\].RFW.CG\[1\]/GCLK DW[14] VGND VGND VPWR VPWR
+ REGF\[14\].RFW.BIT\[14\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[15\].RFW.BIT\[10\].OBUF1 REGF\[15\].RFW.BIT\[10\].FF/Q REGF\[15\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[10] sky130_fd_sc_hd__ebufn_2
XREGF\[30\].RFW.BIT\[17\].FF REGF\[30\].RFW.CG\[2\]/GCLK DW[17] VGND VGND VPWR VPWR
+ REGF\[30\].RFW.BIT\[17\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[31\].RFW.BIT\[1\].OBUF2 REGF\[31\].RFW.BIT\[1\].FF/Q REGF\[31\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[1] sky130_fd_sc_hd__ebufn_2
Xgenblk1.RFW0.BIT\[26\].OBUF1 genblk1.RFW0.TIE\[3\]/LO genblk1.RFW0.INV1\[3\]/Y VGND
+ VGND VPWR VPWR DA[26] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[26\].OBUF2 REGF\[16\].RFW.BIT\[26\].FF/Q REGF\[16\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[26] sky130_fd_sc_hd__ebufn_2
XDEC1.D2.AND0 DEC1.D2.AND7/A DEC1.D2.AND7/B DEC1.D2.AND7/C DEC1.D2.AND7/D VGND VGND
+ VPWR VPWR DEC1.D2.AND0/Y sky130_fd_sc_hd__nor4b_2
Xfill_31_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_24_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_17_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[21\].RFW.BIT\[15\].OBUF2 REGF\[21\].RFW.BIT\[15\].FF/Q REGF\[21\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[15] sky130_fd_sc_hd__ebufn_2
XREGF\[25\].RFW.BIT\[24\].FF REGF\[25\].RFW.CG\[3\]/GCLK DW[24] VGND VGND VPWR VPWR
+ REGF\[25\].RFW.BIT\[24\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[19\].RFW.BIT\[11\].OBUF2 REGF\[19\].RFW.BIT\[11\].FF/Q REGF\[19\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[11] sky130_fd_sc_hd__ebufn_2
XREGF\[11\].RFW.BIT\[13\].OBUF1 REGF\[11\].RFW.BIT\[13\].FF/Q REGF\[11\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[13] sky130_fd_sc_hd__ebufn_2
Xfill_17_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_17_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_17_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_17_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_17_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.BIT\[29\].OBUF2 REGF\[12\].RFW.BIT\[29\].FF/Q REGF\[12\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[29] sky130_fd_sc_hd__ebufn_2
Xfill_33_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_33_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xtap_58_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC0.D3.AND2 DEC0.D3.AND7/C DEC0.D3.AND7/A DEC0.D3.AND7/B DEC0.D3.AND7/D VGND VGND
+ VPWR VPWR DEC0.D3.AND2/X sky130_fd_sc_hd__and4bb_2
Xfill_58_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_58_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_5_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.BIT\[21\].OBUF2 REGF\[3\].RFW.BIT\[21\].FF/Q REGF\[3\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[21] sky130_fd_sc_hd__ebufn_2
Xfill_58_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_5_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_5_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[15\].RFW.BIT\[14\].OBUF2 REGF\[15\].RFW.BIT\[14\].FF/Q REGF\[15\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[14] sky130_fd_sc_hd__ebufn_2
Xfill_10_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[9\].RFW.INV1\[1\] DEC0.D1.AND1/X VGND VGND VPWR VPWR REGF\[9\].RFW.INV1\[1\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_22_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.BIT\[30\].OBUF2 REGF\[12\].RFW.BIT\[30\].FF/Q REGF\[12\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[30] sky130_fd_sc_hd__ebufn_2
XREGF\[11\].RFW.BIT\[17\].OBUF2 REGF\[11\].RFW.BIT\[17\].FF/Q REGF\[11\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[17] sky130_fd_sc_hd__ebufn_2
XREGF\[11\].RFW.BIT\[22\].FF REGF\[11\].RFW.CG\[2\]/GCLK DW[22] VGND VGND VPWR VPWR
+ REGF\[11\].RFW.BIT\[22\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_44_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.CG\[3\] CLK REGF\[6\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[6\].RFW.CG\[3\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_2_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_28_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_28_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_28_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[27\].RFW.BIT\[27\].OBUF1 REGF\[27\].RFW.BIT\[27\].FF/Q REGF\[27\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[27] sky130_fd_sc_hd__ebufn_2
Xfill_44_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_44_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_44_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.CGAND DEC2.D0.AND3/X WE VGND VGND VPWR VPWR REGF\[3\].RFW.CGAND/X sky130_fd_sc_hd__and2_1
Xgenblk1.RFW0.BIT\[31\].OBUF2 genblk1.RFW0.TIE\[7\]/LO genblk1.RFW0.INV2\[3\]/Y VGND
+ VGND VPWR VPWR DB[31] sky130_fd_sc_hd__ebufn_2
Xfill_60_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_60_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_60_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_58_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[5\].RFW.CG\[0\] CLK REGF\[5\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[5\].RFW.CG\[0\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[30\].RFW.BIT\[0\].FF REGF\[30\].RFW.CG\[0\]/GCLK DW[0] VGND VGND VPWR VPWR
+ REGF\[30\].RFW.BIT\[0\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_6_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.BIT\[15\].FF REGF\[6\].RFW.CG\[1\]/GCLK DW[15] VGND VGND VPWR VPWR
+ REGF\[6\].RFW.BIT\[15\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[3\].RFW.INV2\[2\] DEC1.D0.AND3/X VGND VGND VPWR VPWR REGF\[3\].RFW.INV2\[2\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[26\].RFW.BIT\[15\].OBUF1 REGF\[26\].RFW.BIT\[15\].FF/Q REGF\[26\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[15] sky130_fd_sc_hd__ebufn_2
Xfill_14_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_30_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[23\].RFW.INV2\[0\] DEC1.D2.AND7/X VGND VGND VPWR VPWR REGF\[23\].RFW.INV2\[0\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_30_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_30_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[23\].RFW.BIT\[15\].FF REGF\[23\].RFW.CG\[1\]/GCLK DW[15] VGND VGND VPWR VPWR
+ REGF\[23\].RFW.BIT\[15\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_42_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC0.D0.AND5 DEC0.D0.AND7/B DEC0.D0.AND7/A DEC0.D0.AND7/C DEC0.D0.AND7/D VGND VGND
+ VPWR VPWR DEC0.D0.AND5/X sky130_fd_sc_hd__and4b_2
Xtap_35_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_28_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_39_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_39_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_39_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_55_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_55_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_55_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_55_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_2_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[17\].RFW.BIT\[29\].OBUF1 REGF\[17\].RFW.BIT\[29\].FF/Q REGF\[17\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[29] sky130_fd_sc_hd__ebufn_2
Xfill_55_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[22\].RFW.BIT\[18\].OBUF1 REGF\[22\].RFW.BIT\[18\].FF/Q REGF\[22\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[18] sky130_fd_sc_hd__ebufn_2
XREGF\[23\].RFW.BIT\[31\].OBUF1 REGF\[23\].RFW.BIT\[31\].FF/Q REGF\[23\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[31] sky130_fd_sc_hd__ebufn_2
XREGF\[12\].RFW.BIT\[28\].FF REGF\[12\].RFW.CG\[3\]/GCLK DW[28] VGND VGND VPWR VPWR
+ REGF\[12\].RFW.BIT\[28\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[8\].RFW.BIT\[21\].OBUF1 REGF\[8\].RFW.BIT\[21\].FF/Q REGF\[8\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[21] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.BIT\[22\].FF REGF\[18\].RFW.CG\[2\]/GCLK DW[22] VGND VGND VPWR VPWR
+ REGF\[18\].RFW.BIT\[22\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_56_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[13\].RFW.CGAND DEC2.D1.AND5/X WE VGND VGND VPWR VPWR REGF\[13\].RFW.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_49_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_4_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[26\].RFW.BIT\[19\].OBUF2 REGF\[26\].RFW.BIT\[19\].FF/Q REGF\[26\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[19] sky130_fd_sc_hd__ebufn_2
Xtap_14_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[4\].RFW.BIT\[24\].OBUF1 REGF\[4\].RFW.BIT\[24\].FF/Q REGF\[4\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[24] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[17\].OBUF1 REGF\[16\].RFW.BIT\[17\].FF/Q REGF\[16\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[17] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.BIT\[30\].OBUF1 REGF\[17\].RFW.BIT\[30\].FF/Q REGF\[17\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[30] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.INV2\[1\] DEC1.D2.AND2/X VGND VGND VPWR VPWR REGF\[18\].RFW.INV2\[1\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_25_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_25_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_25_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_25_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_25_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_41_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_41_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_41_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_41_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_41_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDEC1.D.AND1 RB[4] RB[3] DEC1.TIE/HI VGND VGND VPWR VPWR DEC1.D.AND1/X sky130_fd_sc_hd__and3b_4
Xtap_40_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.BIT\[23\].FF REGF\[3\].RFW.CG\[2\]/GCLK DW[23] VGND VGND VPWR VPWR
+ REGF\[3\].RFW.BIT\[23\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_33_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.BIT\[10\].FF REGF\[31\].RFW.CG\[1\]/GCLK DW[10] VGND VGND VPWR VPWR
+ REGF\[31\].RFW.BIT\[10\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[8\].RFW.BIT\[25\].OBUF2 REGF\[8\].RFW.BIT\[25\].FF/Q REGF\[8\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[25] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[20\].OBUF2 REGF\[26\].RFW.BIT\[20\].FF/Q REGF\[26\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[20] sky130_fd_sc_hd__ebufn_2
XREGF\[20\].RFW.BIT\[23\].FF REGF\[20\].RFW.CG\[2\]/GCLK DW[23] VGND VGND VPWR VPWR
+ REGF\[20\].RFW.BIT\[23\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_61_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.BIT\[12\].OBUF1 REGF\[3\].RFW.BIT\[12\].FF/Q REGF\[3\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[12] sky130_fd_sc_hd__ebufn_2
Xfill_54_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[14\].RFW.INV1\[2\] DEC0.D1.AND6/X VGND VGND VPWR VPWR REGF\[14\].RFW.INV1\[2\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_47_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_3_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_3_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_2_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XREGF\[4\].RFW.BIT\[28\].OBUF2 REGF\[4\].RFW.BIT\[28\].FF/Q REGF\[4\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[28] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.BIT\[28\].FF REGF\[19\].RFW.CG\[3\]/GCLK DW[28] VGND VGND VPWR VPWR
+ REGF\[19\].RFW.BIT\[28\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_11_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_11_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_11_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[15\].RFW.BIT\[30\].FF REGF\[15\].RFW.CG\[3\]/GCLK DW[30] VGND VGND VPWR VPWR
+ REGF\[15\].RFW.BIT\[30\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[22\].RFW.BIT\[23\].OBUF2 REGF\[22\].RFW.BIT\[23\].FF/Q REGF\[22\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[23] sky130_fd_sc_hd__ebufn_2
Xtap_12_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[7\].RFW.BIT\[13\].OBUF2 REGF\[7\].RFW.BIT\[13\].FF/Q REGF\[7\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[13] sky130_fd_sc_hd__ebufn_2
Xtap_5_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_36_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_36_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_36_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_52_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_52_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[12\].RFW.BIT\[21\].OBUF1 REGF\[12\].RFW.BIT\[21\].FF/Q REGF\[12\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[21] sky130_fd_sc_hd__ebufn_2
Xfill_52_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_8_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_8_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_40_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_26_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_19_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgenblk1.RFW0.BIT\[22\].OBUF1 genblk1.RFW0.TIE\[2\]/LO genblk1.RFW0.INV1\[2\]/Y VGND
+ VGND VPWR VPWR DA[22] sky130_fd_sc_hd__ebufn_2
XREGF\[3\].RFW.BIT\[16\].OBUF2 REGF\[3\].RFW.BIT\[16\].FF/Q REGF\[3\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[16] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[22\].OBUF2 REGF\[16\].RFW.BIT\[22\].FF/Q REGF\[16\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[22] sky130_fd_sc_hd__ebufn_2
XREGF\[10\].RFW.BIT\[19\].FF REGF\[10\].RFW.CG\[2\]/GCLK DW[19] VGND VGND VPWR VPWR
+ REGF\[10\].RFW.BIT\[19\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[4\].RFW.BIT\[29\].FF REGF\[4\].RFW.CG\[3\]/GCLK DW[29] VGND VGND VPWR VPWR
+ REGF\[4\].RFW.BIT\[29\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[21\].RFW.BIT\[11\].OBUF2 REGF\[21\].RFW.BIT\[11\].FF/Q REGF\[21\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[11] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[13\].FF REGF\[16\].RFW.CG\[1\]/GCLK DW[13] VGND VGND VPWR VPWR
+ REGF\[16\].RFW.BIT\[13\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_52_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_22_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_22_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_22_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[21\].RFW.BIT\[29\].FF REGF\[21\].RFW.CG\[3\]/GCLK DW[29] VGND VGND VPWR VPWR
+ REGF\[21\].RFW.BIT\[29\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_10_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.BIT\[25\].OBUF2 REGF\[12\].RFW.BIT\[25\].FF/Q REGF\[12\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[25] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[23\].FF REGF\[27\].RFW.CG\[2\]/GCLK DW[23] VGND VGND VPWR VPWR
+ REGF\[27\].RFW.BIT\[23\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_47_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_47_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_47_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_47_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xtap_3_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_47_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[1\].RFW.INV1\[0\] DEC0.D0.AND1/X VGND VGND VPWR VPWR REGF\[1\].RFW.INV1\[0\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[15\].RFW.BIT\[10\].OBUF2 REGF\[15\].RFW.BIT\[10\].FF/Q REGF\[15\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[10] sky130_fd_sc_hd__ebufn_2
XREGF\[1\].RFW.BIT\[14\].FF REGF\[1\].RFW.CG\[1\]/GCLK DW[14] VGND VGND VPWR VPWR
+ REGF\[1\].RFW.BIT\[14\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xgenblk1.RFW0.BIT\[26\].OBUF2 genblk1.RFW0.TIE\[7\]/LO genblk1.RFW0.INV2\[3\]/Y VGND
+ VGND VPWR VPWR DB[26] sky130_fd_sc_hd__ebufn_2
XDEC1.D2.AND1 DEC1.D2.AND7/C DEC1.D2.AND7/B DEC1.D2.AND7/A DEC1.D2.AND7/D VGND VGND
+ VPWR VPWR DEC1.D2.AND1/X sky130_fd_sc_hd__and4bb_2
Xfill_31_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_24_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_9_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[2\].RFW.CG\[2\] CLK REGF\[2\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[2\].RFW.CG\[2\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[11\].RFW.BIT\[13\].OBUF2 REGF\[11\].RFW.BIT\[13\].FF/Q REGF\[11\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[13] sky130_fd_sc_hd__ebufn_2
Xfill_17_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_17_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[9\].RFW.BIT\[28\].OBUF1 REGF\[9\].RFW.BIT\[28\].FF/Q REGF\[9\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[28] sky130_fd_sc_hd__ebufn_2
Xfill_17_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[2\].RFW.CGAND DEC2.D0.AND2/X WE VGND VGND VPWR VPWR REGF\[2\].RFW.CGAND/X sky130_fd_sc_hd__and2_1
Xfill_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_33_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_33_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[28\].RFW.CG\[1\] CLK REGF\[28\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[28\].RFW.CG\[1\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[27\].RFW.BIT\[23\].OBUF1 REGF\[27\].RFW.BIT\[23\].FF/Q REGF\[27\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[23] sky130_fd_sc_hd__ebufn_2
Xtap_58_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC0.D3.AND3 DEC0.D3.AND7/C DEC0.D3.AND7/B DEC0.D3.AND7/A DEC0.D3.AND7/D VGND VGND
+ VPWR VPWR DEC0.D3.AND3/X sky130_fd_sc_hd__and4b_2
XREGF\[17\].RFW.BIT\[19\].FF REGF\[17\].RFW.CG\[2\]/GCLK DW[19] VGND VGND VPWR VPWR
+ REGF\[17\].RFW.BIT\[19\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_58_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_58_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[7\].RFW.BIT\[31\].FF REGF\[7\].RFW.CG\[3\]/GCLK DW[31] VGND VGND VPWR VPWR
+ REGF\[7\].RFW.BIT\[31\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[13\].RFW.BIT\[21\].FF REGF\[13\].RFW.CG\[2\]/GCLK DW[21] VGND VGND VPWR VPWR
+ REGF\[13\].RFW.BIT\[21\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_58_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_5_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_5_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC1.D2.ABUF\[0\] RB[0] VGND VGND VPWR VPWR DEC1.D2.AND7/A sky130_fd_sc_hd__clkbuf_2
XREGF\[23\].RFW.BIT\[26\].OBUF1 REGF\[23\].RFW.BIT\[26\].FF/Q REGF\[23\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[26] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.BIT\[29\].FF REGF\[28\].RFW.CG\[3\]/GCLK DW[29] VGND VGND VPWR VPWR
+ REGF\[28\].RFW.BIT\[29\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[24\].RFW.BIT\[31\].FF REGF\[24\].RFW.CG\[3\]/GCLK DW[31] VGND VGND VPWR VPWR
+ REGF\[24\].RFW.BIT\[31\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[8\].RFW.BIT\[16\].OBUF1 REGF\[8\].RFW.BIT\[16\].FF/Q REGF\[8\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[16] sky130_fd_sc_hd__ebufn_2
Xfill_22_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_15_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.INV2\[0\] DEC1.D3.AND7/X VGND VGND VPWR VPWR REGF\[31\].RFW.INV2\[0\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[26\].RFW.BIT\[11\].OBUF1 REGF\[26\].RFW.BIT\[11\].FF/Q REGF\[26\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[11] sky130_fd_sc_hd__ebufn_2
Xtap_44_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[8\].RFW.BIT\[14\].FF REGF\[8\].RFW.CG\[1\]/GCLK DW[14] VGND VGND VPWR VPWR
+ REGF\[8\].RFW.BIT\[14\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_28_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[16\].RFW.CG\[1\] CLK REGF\[16\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[16\].RFW.CG\[1\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_28_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_28_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[27\].RFW.BIT\[27\].OBUF2 REGF\[27\].RFW.BIT\[27\].FF/Q REGF\[27\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[27] sky130_fd_sc_hd__ebufn_2
Xfill_44_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_44_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_44_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_60_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[4\].RFW.BIT\[19\].OBUF1 REGF\[4\].RFW.BIT\[19\].FF/Q REGF\[4\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[19] sky130_fd_sc_hd__ebufn_2
Xfill_60_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_60_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[17\].RFW.BIT\[25\].OBUF1 REGF\[17\].RFW.BIT\[25\].FF/Q REGF\[17\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[25] sky130_fd_sc_hd__ebufn_2
XREGF\[22\].RFW.BIT\[14\].OBUF1 REGF\[22\].RFW.BIT\[14\].FF/Q REGF\[22\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[14] sky130_fd_sc_hd__ebufn_2
XREGF\[12\].RFW.CGAND DEC2.D1.AND4/X WE VGND VGND VPWR VPWR REGF\[12\].RFW.CGAND/X
+ sky130_fd_sc_hd__and2_1
XREGF\[25\].RFW.BIT\[14\].FF REGF\[25\].RFW.CG\[1\]/GCLK DW[14] VGND VGND VPWR VPWR
+ REGF\[25\].RFW.BIT\[14\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[6\].RFW.INV2\[3\] DEC1.D0.AND6/X VGND VGND VPWR VPWR REGF\[6\].RFW.INV2\[3\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_6_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[18\].RFW.BIT\[1\].FF REGF\[18\].RFW.CG\[0\]/GCLK DW[1] VGND VGND VPWR VPWR
+ REGF\[18\].RFW.BIT\[1\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[14\].RFW.BIT\[27\].FF REGF\[14\].RFW.CG\[3\]/GCLK DW[27] VGND VGND VPWR VPWR
+ REGF\[14\].RFW.BIT\[27\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[10\].RFW.INV2\[0\] DEC1.D1.AND2/X VGND VGND VPWR VPWR REGF\[10\].RFW.INV2\[0\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[26\].RFW.BIT\[15\].OBUF2 REGF\[26\].RFW.BIT\[15\].FF/Q REGF\[26\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[15] sky130_fd_sc_hd__ebufn_2
XREGF\[13\].RFW.BIT\[28\].OBUF1 REGF\[13\].RFW.BIT\[28\].FF/Q REGF\[13\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[28] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.INV2\[1\] DEC1.D3.AND2/X VGND VGND VPWR VPWR REGF\[26\].RFW.INV2\[1\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_14_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_14_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[17\].RFW.BIT\[3\].FF REGF\[17\].RFW.CG\[0\]/GCLK DW[3] VGND VGND VPWR VPWR
+ REGF\[17\].RFW.BIT\[3\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[4\].RFW.BIT\[20\].OBUF1 REGF\[4\].RFW.BIT\[20\].FF/Q REGF\[4\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[20] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[13\].OBUF1 REGF\[16\].RFW.BIT\[13\].FF/Q REGF\[16\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[13] sky130_fd_sc_hd__ebufn_2
Xfill_30_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_30_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_30_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xtap_42_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC0.D0.AND6 DEC0.D0.AND7/A DEC0.D0.AND7/B DEC0.D0.AND7/C DEC0.D0.AND7/D VGND VGND
+ VPWR VPWR DEC0.D0.AND6/X sky130_fd_sc_hd__and4b_2
Xtap_28_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_39_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[16\].RFW.BIT\[5\].FF REGF\[16\].RFW.CG\[0\]/GCLK DW[5] VGND VGND VPWR VPWR
+ REGF\[16\].RFW.BIT\[5\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_55_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_55_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_55_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_55_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_2_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[17\].RFW.BIT\[29\].OBUF2 REGF\[17\].RFW.BIT\[29\].FF/Q REGF\[17\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[29] sky130_fd_sc_hd__ebufn_2
Xfill_55_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC0.D3.ABUF\[1\] RA[1] VGND VGND VPWR VPWR DEC0.D3.AND7/B sky130_fd_sc_hd__clkbuf_2
XREGF\[22\].RFW.BIT\[18\].OBUF2 REGF\[22\].RFW.BIT\[18\].FF/Q REGF\[22\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[18] sky130_fd_sc_hd__ebufn_2
XREGF\[23\].RFW.BIT\[31\].OBUF2 REGF\[23\].RFW.BIT\[31\].FF/Q REGF\[23\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[31] sky130_fd_sc_hd__ebufn_2
XREGF\[8\].RFW.BIT\[21\].OBUF2 REGF\[8\].RFW.BIT\[21\].FF/Q REGF\[8\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[21] sky130_fd_sc_hd__ebufn_2
XREGF\[15\].RFW.BIT\[7\].FF REGF\[15\].RFW.CG\[0\]/GCLK DW[7] VGND VGND VPWR VPWR
+ REGF\[15\].RFW.BIT\[7\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[22\].RFW.INV1\[2\] DEC0.D2.AND6/X VGND VGND VPWR VPWR REGF\[22\].RFW.INV1\[2\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_56_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[12\].RFW.BIT\[16\].OBUF1 REGF\[12\].RFW.BIT\[16\].FF/Q REGF\[12\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[16] sky130_fd_sc_hd__ebufn_2
Xgenblk1.RFW0.INV1\[0\] DEC0.D0.AND0/Y VGND VGND VPWR VPWR genblk1.RFW0.INV1\[0\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_49_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[5\].RFW.BIT\[22\].FF REGF\[5\].RFW.CG\[2\]/GCLK DW[22] VGND VGND VPWR VPWR
+ REGF\[5\].RFW.BIT\[22\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[11\].RFW.BIT\[12\].FF REGF\[11\].RFW.CG\[1\]/GCLK DW[12] VGND VGND VPWR VPWR
+ REGF\[11\].RFW.BIT\[12\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_4_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[14\].RFW.BIT\[9\].FF REGF\[14\].RFW.CG\[1\]/GCLK DW[9] VGND VGND VPWR VPWR
+ REGF\[14\].RFW.BIT\[9\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xgenblk1.RFW0.BIT\[17\].OBUF1 genblk1.RFW0.TIE\[2\]/LO genblk1.RFW0.INV1\[2\]/Y VGND
+ VGND VPWR VPWR DA[17] sky130_fd_sc_hd__ebufn_2
Xtap_14_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[4\].RFW.BIT\[24\].OBUF2 REGF\[4\].RFW.BIT\[24\].FF/Q REGF\[4\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[24] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.BIT\[5\].FF REGF\[29\].RFW.CG\[0\]/GCLK DW[5] VGND VGND VPWR VPWR
+ REGF\[29\].RFW.BIT\[5\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[16\].RFW.BIT\[17\].OBUF2 REGF\[16\].RFW.BIT\[17\].FF/Q REGF\[16\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[17] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.BIT\[30\].OBUF2 REGF\[17\].RFW.BIT\[30\].FF/Q REGF\[17\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[30] sky130_fd_sc_hd__ebufn_2
XREGF\[22\].RFW.BIT\[22\].FF REGF\[22\].RFW.CG\[2\]/GCLK DW[22] VGND VGND VPWR VPWR
+ REGF\[22\].RFW.BIT\[22\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_25_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_25_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_25_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_25_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_41_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_41_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_41_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[28\].RFW.BIT\[7\].FF REGF\[28\].RFW.CG\[0\]/GCLK DW[7] VGND VGND VPWR VPWR
+ REGF\[28\].RFW.BIT\[7\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_41_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC1.D.AND2 RB[3] RB[4] DEC1.TIE/HI VGND VGND VPWR VPWR DEC1.D.AND2/X sky130_fd_sc_hd__and3b_4
Xtap_40_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[27\].RFW.BIT\[9\].FF REGF\[27\].RFW.CG\[1\]/GCLK DW[9] VGND VGND VPWR VPWR
+ REGF\[27\].RFW.BIT\[9\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_15_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[17\].RFW.INV1\[3\] DEC0.D2.AND1/X VGND VGND VPWR VPWR REGF\[17\].RFW.INV1\[3\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_61_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[3\].RFW.BIT\[12\].OBUF2 REGF\[3\].RFW.BIT\[12\].FF/Q REGF\[3\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[12] sky130_fd_sc_hd__ebufn_2
Xfill_54_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_47_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_3_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_2_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_11_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_11_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_12_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.BIT\[28\].FF REGF\[6\].RFW.CG\[3\]/GCLK DW[28] VGND VGND VPWR VPWR
+ REGF\[6\].RFW.BIT\[28\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[12\].RFW.BIT\[18\].FF REGF\[12\].RFW.CG\[2\]/GCLK DW[18] VGND VGND VPWR VPWR
+ REGF\[12\].RFW.BIT\[18\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[2\].RFW.BIT\[30\].FF REGF\[2\].RFW.CG\[3\]/GCLK DW[30] VGND VGND VPWR VPWR
+ REGF\[2\].RFW.BIT\[30\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_5_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_36_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_36_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_36_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[18\].RFW.BIT\[12\].FF REGF\[18\].RFW.CG\[1\]/GCLK DW[12] VGND VGND VPWR VPWR
+ REGF\[18\].RFW.BIT\[12\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_52_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_52_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_52_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.BIT\[21\].OBUF2 REGF\[12\].RFW.BIT\[21\].FF/Q REGF\[12\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[21] sky130_fd_sc_hd__ebufn_2
Xfill_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_8_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[8\].RFW.INV2\[0\] DEC1.D1.AND0/Y VGND VGND VPWR VPWR REGF\[8\].RFW.INV2\[0\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[23\].RFW.BIT\[28\].FF REGF\[23\].RFW.CG\[3\]/GCLK DW[28] VGND VGND VPWR VPWR
+ REGF\[23\].RFW.BIT\[28\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[27\].RFW.BIT\[18\].OBUF1 REGF\[27\].RFW.BIT\[18\].FF/Q REGF\[27\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[18] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.BIT\[31\].OBUF1 REGF\[28\].RFW.BIT\[31\].FF/Q REGF\[28\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[31] sky130_fd_sc_hd__ebufn_2
Xfill_33_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[25\].RFW.CG\[3\] CLK REGF\[25\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[25\].RFW.CG\[3\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_26_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_19_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[29\].RFW.BIT\[22\].FF REGF\[29\].RFW.CG\[2\]/GCLK DW[22] VGND VGND VPWR VPWR
+ REGF\[29\].RFW.BIT\[22\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xgenblk1.RFW0.BIT\[22\].OBUF2 genblk1.RFW0.TIE\[6\]/LO genblk1.RFW0.INV2\[2\]/Y VGND
+ VGND VPWR VPWR DB[22] sky130_fd_sc_hd__ebufn_2
Xfill_52_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_45_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[1\].RFW.CGAND DEC2.D0.AND1/X WE VGND VGND VPWR VPWR REGF\[1\].RFW.CGAND/X sky130_fd_sc_hd__and2_1
XREGF\[3\].RFW.BIT\[13\].FF REGF\[3\].RFW.CG\[1\]/GCLK DW[13] VGND VGND VPWR VPWR
+ REGF\[3\].RFW.BIT\[13\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_0_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[24\].RFW.CG\[0\] CLK REGF\[24\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[24\].RFW.CG\[0\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XDEC2.D1.AND0 DEC2.D1.AND7/A DEC2.D1.AND7/B DEC2.D1.AND7/C DEC2.D1.AND7/D VGND VGND
+ VPWR VPWR DEC2.D1.AND0/Y sky130_fd_sc_hd__nor4b_2
Xfill_22_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_22_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[4\].RFW.INV1\[1\] DEC0.D0.AND4/X VGND VGND VPWR VPWR REGF\[4\].RFW.INV1\[1\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[9\].RFW.BIT\[24\].OBUF1 REGF\[9\].RFW.BIT\[24\].FF/Q REGF\[9\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[24] sky130_fd_sc_hd__ebufn_2
Xtap_10_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_47_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_47_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_47_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_47_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_47_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[20\].RFW.BIT\[13\].FF REGF\[20\].RFW.CG\[1\]/GCLK DW[13] VGND VGND VPWR VPWR
+ REGF\[20\].RFW.BIT\[13\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[13\].RFW.CG\[3\] CLK REGF\[13\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[13\].RFW.CG\[3\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[1\].RFW.BIT\[9\].OBUF1 REGF\[1\].RFW.BIT\[9\].FF/Q REGF\[1\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[9] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[27\].OBUF1 REGF\[5\].RFW.BIT\[27\].FF/Q REGF\[5\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[27] sky130_fd_sc_hd__ebufn_2
XDEC1.D2.AND2 DEC1.D2.AND7/C DEC1.D2.AND7/A DEC1.D2.AND7/B DEC1.D2.AND7/D VGND VGND
+ VPWR VPWR DEC1.D2.AND2/X sky130_fd_sc_hd__and4bb_2
Xfill_31_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[19\].RFW.BIT\[18\].FF REGF\[19\].RFW.CG\[2\]/GCLK DW[18] VGND VGND VPWR VPWR
+ REGF\[19\].RFW.BIT\[18\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_24_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[9\].RFW.BIT\[30\].FF REGF\[9\].RFW.CG\[3\]/GCLK DW[30] VGND VGND VPWR VPWR
+ REGF\[9\].RFW.BIT\[30\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[15\].RFW.BIT\[20\].FF REGF\[15\].RFW.CG\[2\]/GCLK DW[20] VGND VGND VPWR VPWR
+ REGF\[15\].RFW.BIT\[20\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[12\].RFW.BIT\[0\].FF REGF\[12\].RFW.CG\[0\]/GCLK DW[0] VGND VGND VPWR VPWR
+ REGF\[12\].RFW.BIT\[0\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_17_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.BIT\[23\].FF REGF\[31\].RFW.CG\[2\]/GCLK DW[23] VGND VGND VPWR VPWR
+ REGF\[31\].RFW.BIT\[23\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[23\].RFW.BIT\[22\].OBUF1 REGF\[23\].RFW.BIT\[22\].FF/Q REGF\[23\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[22] sky130_fd_sc_hd__ebufn_2
XREGF\[8\].RFW.BIT\[12\].OBUF1 REGF\[8\].RFW.BIT\[12\].FF/Q REGF\[8\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[12] sky130_fd_sc_hd__ebufn_2
Xfill_9_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_9_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.CG\[0\] CLK REGF\[12\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[12\].RFW.CG\[0\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[11\].RFW.BIT\[2\].FF REGF\[11\].RFW.CG\[0\]/GCLK DW[2] VGND VGND VPWR VPWR
+ REGF\[11\].RFW.BIT\[2\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_17_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_17_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_17_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[9\].RFW.BIT\[28\].OBUF2 REGF\[9\].RFW.BIT\[28\].FF/Q REGF\[9\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[28] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[30\].FF REGF\[26\].RFW.CG\[3\]/GCLK DW[30] VGND VGND VPWR VPWR
+ REGF\[26\].RFW.BIT\[30\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_33_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_33_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.BIT\[9\].OBUF1 REGF\[3\].RFW.BIT\[9\].FF/Q REGF\[3\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[9] sky130_fd_sc_hd__ebufn_2
Xtap_58_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC0.D3.AND4 DEC0.D3.AND7/A DEC0.D3.AND7/B DEC0.D3.AND7/C DEC0.D3.AND7/D VGND VGND
+ VPWR VPWR DEC0.D3.AND4/X sky130_fd_sc_hd__and4bb_2
XREGF\[27\].RFW.BIT\[23\].OBUF2 REGF\[27\].RFW.BIT\[23\].FF/Q REGF\[27\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[23] sky130_fd_sc_hd__ebufn_2
XREGF\[10\].RFW.BIT\[4\].FF REGF\[10\].RFW.CG\[0\]/GCLK DW[4] VGND VGND VPWR VPWR
+ REGF\[10\].RFW.BIT\[4\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[11\].RFW.CGAND DEC2.D1.AND3/X WE VGND VGND VPWR VPWR REGF\[11\].RFW.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_58_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_58_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_58_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_5_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[4\].RFW.BIT\[15\].OBUF1 REGF\[4\].RFW.BIT\[15\].FF/Q REGF\[4\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[15] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.BIT\[21\].OBUF1 REGF\[17\].RFW.BIT\[21\].FF/Q REGF\[17\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[21] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.INV1\[0\] DEC0.D2.AND3/X VGND VGND VPWR VPWR REGF\[19\].RFW.INV1\[0\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[4\].RFW.BIT\[19\].FF REGF\[4\].RFW.CG\[2\]/GCLK DW[19] VGND VGND VPWR VPWR
+ REGF\[4\].RFW.BIT\[19\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[25\].RFW.BIT\[0\].FF REGF\[25\].RFW.CG\[0\]/GCLK DW[0] VGND VGND VPWR VPWR
+ REGF\[25\].RFW.BIT\[0\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[22\].RFW.BIT\[10\].OBUF1 REGF\[22\].RFW.BIT\[10\].FF/Q REGF\[22\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[10] sky130_fd_sc_hd__ebufn_2
Xfill_23_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[23\].RFW.BIT\[26\].OBUF2 REGF\[23\].RFW.BIT\[26\].FF/Q REGF\[23\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[26] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[2\].FF REGF\[24\].RFW.CG\[0\]/GCLK DW[2] VGND VGND VPWR VPWR
+ REGF\[24\].RFW.BIT\[2\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[8\].RFW.BIT\[16\].OBUF2 REGF\[8\].RFW.BIT\[16\].FF/Q REGF\[8\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[16] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[9\].OBUF1 REGF\[5\].RFW.BIT\[9\].FF/Q REGF\[5\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[9] sky130_fd_sc_hd__ebufn_2
Xfill_22_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XREGF\[21\].RFW.BIT\[19\].FF REGF\[21\].RFW.CG\[2\]/GCLK DW[19] VGND VGND VPWR VPWR
+ REGF\[21\].RFW.BIT\[19\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_15_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XREGF\[1\].RFW.BIT\[31\].OBUF1 REGF\[1\].RFW.BIT\[31\].FF/Q REGF\[1\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[31] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[13\].FF REGF\[27\].RFW.CG\[1\]/GCLK DW[13] VGND VGND VPWR VPWR
+ REGF\[27\].RFW.BIT\[13\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[13\].RFW.BIT\[24\].OBUF1 REGF\[13\].RFW.BIT\[24\].FF/Q REGF\[13\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[24] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[11\].OBUF2 REGF\[26\].RFW.BIT\[11\].FF/Q REGF\[26\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[11] sky130_fd_sc_hd__ebufn_2
XREGF\[23\].RFW.BIT\[4\].FF REGF\[23\].RFW.CG\[0\]/GCLK DW[4] VGND VGND VPWR VPWR
+ REGF\[23\].RFW.BIT\[4\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_44_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_2_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_28_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_28_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_28_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XREGF\[16\].RFW.BIT\[26\].FF REGF\[16\].RFW.CG\[3\]/GCLK DW[26] VGND VGND VPWR VPWR
+ REGF\[16\].RFW.BIT\[26\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[22\].RFW.BIT\[6\].FF REGF\[22\].RFW.CG\[0\]/GCLK DW[6] VGND VGND VPWR VPWR
+ REGF\[22\].RFW.BIT\[6\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_44_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_44_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_44_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_60_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[4\].RFW.BIT\[19\].OBUF2 REGF\[4\].RFW.BIT\[19\].FF/Q REGF\[4\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[19] sky130_fd_sc_hd__ebufn_2
Xfill_60_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_60_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[30\].RFW.INV1\[2\] DEC0.D3.AND6/X VGND VGND VPWR VPWR REGF\[30\].RFW.INV1\[2\]/Y
+ sky130_fd_sc_hd__inv_4
Xtap_56_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[17\].RFW.BIT\[25\].OBUF2 REGF\[17\].RFW.BIT\[25\].FF/Q REGF\[17\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[25] sky130_fd_sc_hd__ebufn_2
XREGF\[8\].RFW.BIT\[1\].FF REGF\[8\].RFW.CG\[0\]/GCLK DW[1] VGND VGND VPWR VPWR REGF\[8\].RFW.BIT\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[7\].RFW.BIT\[9\].OBUF1 REGF\[7\].RFW.BIT\[9\].FF/Q REGF\[7\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[9] sky130_fd_sc_hd__ebufn_2
XREGF\[22\].RFW.BIT\[14\].OBUF2 REGF\[22\].RFW.BIT\[14\].FF/Q REGF\[22\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[14] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.BIT\[8\].FF REGF\[21\].RFW.CG\[1\]/GCLK DW[8] VGND VGND VPWR VPWR
+ REGF\[21\].RFW.BIT\[8\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[10\].RFW.BIT\[8\].OBUF1 REGF\[10\].RFW.BIT\[8\].FF/Q REGF\[10\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[8] sky130_fd_sc_hd__ebufn_2
XREGF\[13\].RFW.INV2\[1\] DEC1.D1.AND5/X VGND VGND VPWR VPWR REGF\[13\].RFW.INV2\[1\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[7\].RFW.BIT\[3\].FF REGF\[7\].RFW.CG\[0\]/GCLK DW[3] VGND VGND VPWR VPWR REGF\[7\].RFW.BIT\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[12\].RFW.BIT\[12\].OBUF1 REGF\[12\].RFW.BIT\[12\].FF/Q REGF\[12\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[12] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.INV2\[2\] DEC1.D3.AND5/X VGND VGND VPWR VPWR REGF\[29\].RFW.INV2\[2\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[13\].RFW.BIT\[28\].OBUF2 REGF\[13\].RFW.BIT\[28\].FF/Q REGF\[13\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[28] sky130_fd_sc_hd__ebufn_2
XREGF\[6\].RFW.BIT\[5\].FF REGF\[6\].RFW.CG\[0\]/GCLK DW[5] VGND VGND VPWR VPWR REGF\[6\].RFW.BIT\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[1\].RFW.BIT\[27\].FF REGF\[1\].RFW.CG\[3\]/GCLK DW[27] VGND VGND VPWR VPWR
+ REGF\[1\].RFW.BIT\[27\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_14_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[9\].RFW.BIT\[9\].OBUF1 REGF\[9\].RFW.BIT\[9\].FF/Q REGF\[9\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[9] sky130_fd_sc_hd__ebufn_2
XREGF\[7\].RFW.BIT\[21\].FF REGF\[7\].RFW.CG\[2\]/GCLK DW[21] VGND VGND VPWR VPWR
+ REGF\[7\].RFW.BIT\[21\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[4\].RFW.BIT\[20\].OBUF2 REGF\[4\].RFW.BIT\[20\].FF/Q REGF\[4\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[20] sky130_fd_sc_hd__ebufn_2
XREGF\[13\].RFW.BIT\[11\].FF REGF\[13\].RFW.CG\[1\]/GCLK DW[11] VGND VGND VPWR VPWR
+ REGF\[13\].RFW.BIT\[11\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xgenblk1.RFW0.BIT\[13\].OBUF1 genblk1.RFW0.TIE\[1\]/LO genblk1.RFW0.INV1\[1\]/Y VGND
+ VGND VPWR VPWR DA[13] sky130_fd_sc_hd__ebufn_2
Xfill_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[16\].RFW.BIT\[13\].OBUF2 REGF\[16\].RFW.BIT\[13\].FF/Q REGF\[16\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[13] sky130_fd_sc_hd__ebufn_2
Xfill_30_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_30_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC0.D0.AND7 DEC0.D0.AND7/A DEC0.D0.AND7/B DEC0.D0.AND7/C DEC0.D0.AND7/D VGND VGND
+ VPWR VPWR DEC0.D0.AND7/X sky130_fd_sc_hd__and4_2
Xtap_42_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.BIT\[8\].OBUF1 REGF\[12\].RFW.BIT\[8\].FF/Q REGF\[12\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[8] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[7\].FF REGF\[5\].RFW.CG\[0\]/GCLK DW[7] VGND VGND VPWR VPWR REGF\[5\].RFW.BIT\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xtap_28_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_39_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_39_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_55_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_55_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_55_14 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_55_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_55_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[25\].RFW.INV1\[3\] DEC0.D3.AND1/X VGND VGND VPWR VPWR REGF\[25\].RFW.INV1\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[2\].RFW.BIT\[7\].OBUF1 REGF\[2\].RFW.BIT\[7\].FF/Q REGF\[2\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[7] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.BIT\[19\].FF REGF\[28\].RFW.CG\[2\]/GCLK DW[19] VGND VGND VPWR VPWR
+ REGF\[28\].RFW.BIT\[19\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[24\].RFW.BIT\[21\].FF REGF\[24\].RFW.CG\[2\]/GCLK DW[21] VGND VGND VPWR VPWR
+ REGF\[24\].RFW.BIT\[21\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[4\].RFW.BIT\[9\].FF REGF\[4\].RFW.CG\[1\]/GCLK DW[9] VGND VGND VPWR VPWR REGF\[4\].RFW.BIT\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xfill_56_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.BIT\[16\].OBUF2 REGF\[12\].RFW.BIT\[16\].FF/Q REGF\[12\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[16] sky130_fd_sc_hd__ebufn_2
Xfill_49_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_4_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[14\].RFW.BIT\[8\].OBUF1 REGF\[14\].RFW.BIT\[8\].FF/Q REGF\[14\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[8] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.BIT\[26\].OBUF1 REGF\[28\].RFW.BIT\[26\].FF/Q REGF\[28\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[26] sky130_fd_sc_hd__ebufn_2
XDEC0.D1.ABUF\[0\] RA[0] VGND VGND VPWR VPWR DEC0.D1.AND7/A sky130_fd_sc_hd__clkbuf_2
Xgenblk1.RFW0.BIT\[17\].OBUF2 genblk1.RFW0.TIE\[6\]/LO genblk1.RFW0.INV2\[2\]/Y VGND
+ VGND VPWR VPWR DB[17] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.BIT\[7\].OBUF1 REGF\[4\].RFW.BIT\[7\].FF/Q REGF\[4\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[7] sky130_fd_sc_hd__ebufn_2
Xfill_25_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_25_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xtap_8_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_25_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_41_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_41_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_41_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC1.D.AND3 RB[4] RB[3] DEC1.TIE/HI VGND VGND VPWR VPWR DEC1.D.AND3/X sky130_fd_sc_hd__and3_4
Xtap_40_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_33_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[21\].RFW.CG\[2\] CLK REGF\[21\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[21\].RFW.CG\[2\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[24\].RFW.BIT\[29\].OBUF1 REGF\[24\].RFW.BIT\[29\].FF/Q REGF\[24\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[29] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[8\].OBUF1 REGF\[16\].RFW.BIT\[8\].FF/Q REGF\[16\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[8] sky130_fd_sc_hd__ebufn_2
XREGF\[30\].RFW.BIT\[31\].OBUF1 REGF\[30\].RFW.BIT\[31\].FF/Q REGF\[30\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[31] sky130_fd_sc_hd__ebufn_2
XREGF\[9\].RFW.BIT\[19\].OBUF1 REGF\[9\].RFW.BIT\[19\].FF/Q REGF\[9\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[19] sky130_fd_sc_hd__ebufn_2
XREGF\[8\].RFW.BIT\[27\].FF REGF\[8\].RFW.CG\[3\]/GCLK DW[27] VGND VGND VPWR VPWR
+ REGF\[8\].RFW.BIT\[27\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[14\].RFW.BIT\[17\].FF REGF\[14\].RFW.CG\[2\]/GCLK DW[17] VGND VGND VPWR VPWR
+ REGF\[14\].RFW.BIT\[17\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_15_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_15_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[27\].RFW.BIT\[14\].OBUF1 REGF\[27\].RFW.BIT\[14\].FF/Q REGF\[27\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[14] sky130_fd_sc_hd__ebufn_2
Xfill_31_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.BIT\[7\].OBUF1 REGF\[6\].RFW.BIT\[7\].FF/Q REGF\[6\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[7] sky130_fd_sc_hd__ebufn_2
Xfill_61_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_54_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_47_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_2_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[25\].RFW.BIT\[27\].FF REGF\[25\].RFW.CG\[3\]/GCLK DW[27] VGND VGND VPWR VPWR
+ REGF\[25\].RFW.BIT\[27\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_11_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.BIT\[28\].OBUF1 REGF\[18\].RFW.BIT\[28\].FF/Q REGF\[18\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[28] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.BIT\[8\].OBUF1 REGF\[18\].RFW.BIT\[8\].FF/Q REGF\[18\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[8] sky130_fd_sc_hd__ebufn_2
Xtap_12_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[23\].RFW.BIT\[17\].OBUF1 REGF\[23\].RFW.BIT\[17\].FF/Q REGF\[23\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[17] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[30\].OBUF1 REGF\[24\].RFW.BIT\[30\].FF/Q REGF\[24\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[30] sky130_fd_sc_hd__ebufn_2
Xfill_36_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_36_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_36_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[9\].RFW.BIT\[20\].OBUF1 REGF\[9\].RFW.BIT\[20\].FF/Q REGF\[9\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[20] sky130_fd_sc_hd__ebufn_2
XREGF\[8\].RFW.BIT\[7\].OBUF1 REGF\[8\].RFW.BIT\[7\].FF/Q REGF\[8\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[7] sky130_fd_sc_hd__ebufn_2
Xfill_52_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_52_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_52_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[5\].RFW.BIT\[12\].FF REGF\[5\].RFW.CG\[1\]/GCLK DW[12] VGND VGND VPWR VPWR
+ REGF\[5\].RFW.BIT\[12\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_8_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[11\].RFW.BIT\[6\].OBUF1 REGF\[11\].RFW.BIT\[6\].FF/Q REGF\[11\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[6] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[18\].OBUF2 REGF\[27\].RFW.BIT\[18\].FF/Q REGF\[27\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[18] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.BIT\[31\].OBUF2 REGF\[28\].RFW.BIT\[31\].FF/Q REGF\[28\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[31] sky130_fd_sc_hd__ebufn_2
Xfill_26_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[1\].RFW.BIT\[5\].OBUF1 REGF\[1\].RFW.BIT\[5\].FF/Q REGF\[1\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[5] sky130_fd_sc_hd__ebufn_2
Xfill_19_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[5\].RFW.BIT\[23\].OBUF1 REGF\[5\].RFW.BIT\[23\].FF/Q REGF\[5\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[23] sky130_fd_sc_hd__ebufn_2
XREGF\[22\].RFW.BIT\[12\].FF REGF\[22\].RFW.CG\[1\]/GCLK DW[12] VGND VGND VPWR VPWR
+ REGF\[22\].RFW.BIT\[12\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[17\].RFW.BIT\[16\].OBUF1 REGF\[17\].RFW.BIT\[16\].FF/Q REGF\[17\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[16] sky130_fd_sc_hd__ebufn_2
Xfill_52_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[7\].RFW.INV1\[2\] DEC0.D0.AND7/X VGND VGND VPWR VPWR REGF\[7\].RFW.INV1\[2\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_45_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_38_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XREGF\[13\].RFW.BIT\[6\].OBUF1 REGF\[13\].RFW.BIT\[6\].FF/Q REGF\[13\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[6] sky130_fd_sc_hd__ebufn_2
XREGF\[11\].RFW.BIT\[25\].FF REGF\[11\].RFW.CG\[3\]/GCLK DW[25] VGND VGND VPWR VPWR
+ REGF\[11\].RFW.BIT\[25\].FF/Q sky130_fd_sc_hd__dfxtp_1
XDEC2.D1.AND1 DEC2.D1.AND7/C DEC2.D1.AND7/B DEC2.D1.AND7/A DEC2.D1.AND7/D VGND VGND
+ VPWR VPWR DEC2.D1.AND1/X sky130_fd_sc_hd__and4bb_2
Xfill_22_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[9\].RFW.BIT\[24\].OBUF2 REGF\[9\].RFW.BIT\[24\].FF/Q REGF\[9\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[24] sky130_fd_sc_hd__ebufn_2
XREGF\[10\].RFW.CGAND DEC2.D1.AND2/X WE VGND VGND VPWR VPWR REGF\[10\].RFW.CGAND/X
+ sky130_fd_sc_hd__and2_1
XREGF\[27\].RFW.INV1\[0\] DEC0.D3.AND3/X VGND VGND VPWR VPWR REGF\[27\].RFW.INV1\[0\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[1\].RFW.BIT\[26\].OBUF1 REGF\[1\].RFW.BIT\[26\].FF/Q REGF\[1\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[26] sky130_fd_sc_hd__ebufn_2
Xtap_10_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.BIT\[5\].OBUF1 REGF\[3\].RFW.BIT\[5\].FF/Q REGF\[3\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[5] sky130_fd_sc_hd__ebufn_2
XREGF\[13\].RFW.BIT\[19\].OBUF1 REGF\[13\].RFW.BIT\[19\].FF/Q REGF\[13\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[19] sky130_fd_sc_hd__ebufn_2
Xfill_47_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_47_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_47_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_47_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_47_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[2\].RFW.BIT\[0\].FF REGF\[2\].RFW.CG\[0\]/GCLK DW[0] VGND VGND VPWR VPWR REGF\[2\].RFW.BIT\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[31\].RFW.BIT\[1\].FF REGF\[31\].RFW.CG\[0\]/GCLK DW[1] VGND VGND VPWR VPWR
+ REGF\[31\].RFW.BIT\[1\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[4\].RFW.BIT\[11\].OBUF1 REGF\[4\].RFW.BIT\[11\].FF/Q REGF\[4\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[11] sky130_fd_sc_hd__ebufn_2
XREGF\[1\].RFW.BIT\[9\].OBUF2 REGF\[1\].RFW.BIT\[9\].FF/Q REGF\[1\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[9] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.CGAND DEC2.D3.AND5/X WE VGND VGND VPWR VPWR REGF\[29\].RFW.CGAND/X
+ sky130_fd_sc_hd__and2_1
XREGF\[5\].RFW.BIT\[27\].OBUF2 REGF\[5\].RFW.BIT\[27\].FF/Q REGF\[5\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[27] sky130_fd_sc_hd__ebufn_2
XDEC1.D2.AND3 DEC1.D2.AND7/C DEC1.D2.AND7/B DEC1.D2.AND7/A DEC1.D2.AND7/D VGND VGND
+ VPWR VPWR DEC1.D2.AND3/X sky130_fd_sc_hd__and4b_2
XREGF\[1\].RFW.BIT\[2\].FF REGF\[1\].RFW.CG\[0\]/GCLK DW[2] VGND VGND VPWR VPWR REGF\[1\].RFW.BIT\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[15\].RFW.BIT\[6\].OBUF1 REGF\[15\].RFW.BIT\[6\].FF/Q REGF\[15\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[6] sky130_fd_sc_hd__ebufn_2
Xfill_31_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[30\].RFW.BIT\[3\].FF REGF\[30\].RFW.CG\[0\]/GCLK DW[3] VGND VGND VPWR VPWR
+ REGF\[30\].RFW.BIT\[3\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_24_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_17_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[23\].RFW.BIT\[22\].OBUF2 REGF\[23\].RFW.BIT\[22\].FF/Q REGF\[23\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[22] sky130_fd_sc_hd__ebufn_2
XREGF\[6\].RFW.BIT\[18\].FF REGF\[6\].RFW.CG\[2\]/GCLK DW[18] VGND VGND VPWR VPWR
+ REGF\[6\].RFW.BIT\[18\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[5\].RFW.BIT\[5\].OBUF1 REGF\[5\].RFW.BIT\[5\].FF/Q REGF\[5\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[5] sky130_fd_sc_hd__ebufn_2
XREGF\[8\].RFW.BIT\[12\].OBUF2 REGF\[8\].RFW.BIT\[12\].FF/Q REGF\[8\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[12] sky130_fd_sc_hd__ebufn_2
Xfill_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_9_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[2\].RFW.BIT\[20\].FF REGF\[2\].RFW.CG\[2\]/GCLK DW[20] VGND VGND VPWR VPWR
+ REGF\[2\].RFW.BIT\[20\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XREGF\[13\].RFW.BIT\[20\].OBUF1 REGF\[13\].RFW.BIT\[20\].FF/Q REGF\[13\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[20] sky130_fd_sc_hd__ebufn_2
XREGF\[1\].RFW.INV2\[3\] DEC1.D0.AND1/X VGND VGND VPWR VPWR REGF\[1\].RFW.INV2\[3\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_17_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_17_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XREGF\[3\].RFW.BIT\[9\].OBUF2 REGF\[3\].RFW.BIT\[9\].FF/Q REGF\[3\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[9] sky130_fd_sc_hd__ebufn_2
Xtap_10_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[23\].RFW.BIT\[18\].FF REGF\[23\].RFW.CG\[2\]/GCLK DW[18] VGND VGND VPWR VPWR
+ REGF\[23\].RFW.BIT\[18\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_58_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC0.D3.AND5 DEC0.D3.AND7/B DEC0.D3.AND7/A DEC0.D3.AND7/C DEC0.D3.AND7/D VGND VGND
+ VPWR VPWR DEC0.D3.AND5/X sky130_fd_sc_hd__and4b_2
XREGF\[17\].RFW.BIT\[6\].OBUF1 REGF\[17\].RFW.BIT\[6\].FF/Q REGF\[17\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[6] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.BIT\[12\].FF REGF\[29\].RFW.CG\[1\]/GCLK DW[12] VGND VGND VPWR VPWR
+ REGF\[29\].RFW.BIT\[12\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_58_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_58_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_58_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[21\].RFW.INV2\[1\] DEC1.D2.AND5/X VGND VGND VPWR VPWR REGF\[21\].RFW.INV2\[1\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[4\].RFW.BIT\[15\].OBUF2 REGF\[4\].RFW.BIT\[15\].FF/Q REGF\[4\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[15] sky130_fd_sc_hd__ebufn_2
Xtap_1_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[17\].RFW.BIT\[21\].OBUF2 REGF\[17\].RFW.BIT\[21\].FF/Q REGF\[17\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[21] sky130_fd_sc_hd__ebufn_2
XREGF\[7\].RFW.BIT\[5\].OBUF1 REGF\[7\].RFW.BIT\[5\].FF/Q REGF\[7\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[5] sky130_fd_sc_hd__ebufn_2
XREGF\[22\].RFW.BIT\[10\].OBUF2 REGF\[22\].RFW.BIT\[10\].FF/Q REGF\[22\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[10] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.BIT\[25\].FF REGF\[18\].RFW.CG\[3\]/GCLK DW[25] VGND VGND VPWR VPWR
+ REGF\[18\].RFW.BIT\[25\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_23_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_23_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[10\].RFW.BIT\[4\].OBUF1 REGF\[10\].RFW.BIT\[4\].FF/Q REGF\[10\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[4] sky130_fd_sc_hd__ebufn_2
XREGF\[30\].RFW.BIT\[30\].FF REGF\[30\].RFW.CG\[3\]/GCLK DW[30] VGND VGND VPWR VPWR
+ REGF\[30\].RFW.BIT\[30\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[5\].RFW.BIT\[9\].OBUF2 REGF\[5\].RFW.BIT\[9\].FF/Q REGF\[5\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[9] sky130_fd_sc_hd__ebufn_2
Xfill_22_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_15_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[1\].RFW.BIT\[31\].OBUF2 REGF\[1\].RFW.BIT\[31\].FF/Q REGF\[1\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[31] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.BIT\[6\].OBUF1 REGF\[19\].RFW.BIT\[6\].FF/Q REGF\[19\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[6] sky130_fd_sc_hd__ebufn_2
XREGF\[13\].RFW.BIT\[24\].OBUF2 REGF\[13\].RFW.BIT\[24\].FF/Q REGF\[13\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[24] sky130_fd_sc_hd__ebufn_2
Xtap_2_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[9\].RFW.BIT\[5\].OBUF1 REGF\[9\].RFW.BIT\[5\].FF/Q REGF\[9\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[5] sky130_fd_sc_hd__ebufn_2
Xfill_28_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_28_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_44_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_44_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.BIT\[4\].OBUF1 REGF\[12\].RFW.BIT\[4\].FF/Q REGF\[12\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[4] sky130_fd_sc_hd__ebufn_2
Xfill_44_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_60_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_60_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_60_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_56_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.BIT\[26\].FF REGF\[3\].RFW.CG\[3\]/GCLK DW[26] VGND VGND VPWR VPWR
+ REGF\[3\].RFW.BIT\[26\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[16\].RFW.INV2\[2\] DEC1.D2.AND0/Y VGND VGND VPWR VPWR REGF\[16\].RFW.INV2\[2\]/Y
+ sky130_fd_sc_hd__inv_4
Xtap_49_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[9\].RFW.BIT\[20\].FF REGF\[9\].RFW.CG\[2\]/GCLK DW[20] VGND VGND VPWR VPWR
+ REGF\[9\].RFW.BIT\[20\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[7\].RFW.BIT\[9\].OBUF2 REGF\[7\].RFW.BIT\[9\].FF/Q REGF\[7\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[9] sky130_fd_sc_hd__ebufn_2
XREGF\[15\].RFW.BIT\[10\].FF REGF\[15\].RFW.CG\[1\]/GCLK DW[10] VGND VGND VPWR VPWR
+ REGF\[15\].RFW.BIT\[10\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[2\].RFW.BIT\[3\].OBUF1 REGF\[2\].RFW.BIT\[3\].FF/Q REGF\[2\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[3] sky130_fd_sc_hd__ebufn_2
XREGF\[31\].RFW.BIT\[13\].FF REGF\[31\].RFW.CG\[1\]/GCLK DW[13] VGND VGND VPWR VPWR
+ REGF\[31\].RFW.BIT\[13\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[10\].RFW.BIT\[8\].OBUF2 REGF\[10\].RFW.BIT\[8\].FF/Q REGF\[10\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[8] sky130_fd_sc_hd__ebufn_2
XREGF\[12\].RFW.BIT\[12\].OBUF2 REGF\[12\].RFW.BIT\[12\].FF/Q REGF\[12\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[12] sky130_fd_sc_hd__ebufn_2
XREGF\[20\].RFW.BIT\[26\].FF REGF\[20\].RFW.CG\[3\]/GCLK DW[26] VGND VGND VPWR VPWR
+ REGF\[20\].RFW.BIT\[26\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[30\].RFW.BIT\[26\].OBUF1 REGF\[30\].RFW.BIT\[26\].FF/Q REGF\[30\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[26] sky130_fd_sc_hd__ebufn_2
Xfill_6_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[26\].RFW.BIT\[20\].FF REGF\[26\].RFW.CG\[2\]/GCLK DW[20] VGND VGND VPWR VPWR
+ REGF\[26\].RFW.BIT\[20\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[14\].RFW.BIT\[4\].OBUF1 REGF\[14\].RFW.BIT\[4\].FF/Q REGF\[14\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[4] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.BIT\[22\].OBUF1 REGF\[28\].RFW.BIT\[22\].FF/Q REGF\[28\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[22] sky130_fd_sc_hd__ebufn_2
Xfill_20_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_14_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.INV1\[3\] DEC0.D1.AND4/X VGND VGND VPWR VPWR REGF\[12\].RFW.INV1\[3\]/Y
+ sky130_fd_sc_hd__inv_4
Xgenblk1.RFW0.BIT\[13\].OBUF2 genblk1.RFW0.TIE\[5\]/LO genblk1.RFW0.INV2\[1\]/Y VGND
+ VGND VPWR VPWR DB[13] sky130_fd_sc_hd__ebufn_2
XREGF\[9\].RFW.BIT\[9\].OBUF2 REGF\[9\].RFW.BIT\[9\].FF/Q REGF\[9\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[9] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.BIT\[3\].OBUF1 REGF\[4\].RFW.BIT\[3\].FF/Q REGF\[4\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[3] sky130_fd_sc_hd__ebufn_2
Xfill_30_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xtap_42_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.BIT\[8\].OBUF2 REGF\[12\].RFW.BIT\[8\].FF/Q REGF\[12\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[8] sky130_fd_sc_hd__ebufn_2
XREGF\[6\].RFW.CG\[1\] CLK REGF\[6\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[6\].RFW.CG\[1\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xtap_28_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_39_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_55_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_55_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_55_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_55_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_55_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[2\].RFW.BIT\[7\].OBUF2 REGF\[2\].RFW.BIT\[7\].FF/Q REGF\[2\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[7] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[25\].OBUF1 REGF\[24\].RFW.BIT\[25\].FF/Q REGF\[24\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[25] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[4\].OBUF1 REGF\[16\].RFW.BIT\[4\].FF/Q REGF\[16\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[4] sky130_fd_sc_hd__ebufn_2
XREGF\[9\].RFW.BIT\[15\].OBUF1 REGF\[9\].RFW.BIT\[15\].FF/Q REGF\[9\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[15] sky130_fd_sc_hd__ebufn_2
Xfill_56_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_29_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[27\].RFW.BIT\[10\].OBUF1 REGF\[27\].RFW.BIT\[10\].FF/Q REGF\[27\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[10] sky130_fd_sc_hd__ebufn_2
Xfill_49_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.BIT\[3\].OBUF1 REGF\[6\].RFW.BIT\[3\].FF/Q REGF\[6\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[3] sky130_fd_sc_hd__ebufn_2
Xfill_4_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[14\].RFW.BIT\[8\].OBUF2 REGF\[14\].RFW.BIT\[8\].FF/Q REGF\[14\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[8] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.BIT\[26\].OBUF2 REGF\[28\].RFW.BIT\[26\].FF/Q REGF\[28\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[26] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[16\].FF REGF\[16\].RFW.CG\[2\]/GCLK DW[16] VGND VGND VPWR VPWR
+ REGF\[16\].RFW.BIT\[16\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[20\].RFW.BIT\[28\].OBUF1 REGF\[20\].RFW.BIT\[28\].FF/Q REGF\[20\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[28] sky130_fd_sc_hd__ebufn_2
XREGF\[3\].RFW.INV2\[0\] DEC1.D0.AND3/X VGND VGND VPWR VPWR REGF\[3\].RFW.INV2\[0\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[5\].RFW.BIT\[18\].OBUF1 REGF\[5\].RFW.BIT\[18\].FF/Q REGF\[5\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[18] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.BIT\[7\].OBUF2 REGF\[4\].RFW.BIT\[7\].FF/Q REGF\[4\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[7] sky130_fd_sc_hd__ebufn_2
XREGF\[6\].RFW.BIT\[31\].OBUF1 REGF\[6\].RFW.BIT\[31\].FF/Q REGF\[6\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[31] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.BIT\[24\].OBUF1 REGF\[18\].RFW.BIT\[24\].FF/Q REGF\[18\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[24] sky130_fd_sc_hd__ebufn_2
Xfill_25_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_8_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.BIT\[4\].OBUF1 REGF\[18\].RFW.BIT\[4\].FF/Q REGF\[18\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[4] sky130_fd_sc_hd__ebufn_2
Xfill_25_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[23\].RFW.BIT\[13\].OBUF1 REGF\[23\].RFW.BIT\[13\].FF/Q REGF\[23\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[13] sky130_fd_sc_hd__ebufn_2
Xfill_41_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_41_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_41_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xtap_40_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[27\].RFW.BIT\[26\].FF REGF\[27\].RFW.CG\[3\]/GCLK DW[26] VGND VGND VPWR VPWR
+ REGF\[27\].RFW.BIT\[26\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_33_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[8\].RFW.BIT\[3\].OBUF1 REGF\[8\].RFW.BIT\[3\].FF/Q REGF\[8\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[3] sky130_fd_sc_hd__ebufn_2
Xgenblk1.RFW0.INV2\[3\] DEC1.D0.AND0/Y VGND VGND VPWR VPWR genblk1.RFW0.INV2\[3\]/Y
+ sky130_fd_sc_hd__inv_4
Xtap_26_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[24\].RFW.BIT\[29\].OBUF2 REGF\[24\].RFW.BIT\[29\].FF/Q REGF\[24\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[29] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[8\].OBUF2 REGF\[16\].RFW.BIT\[8\].FF/Q REGF\[16\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[8] sky130_fd_sc_hd__ebufn_2
XREGF\[30\].RFW.BIT\[31\].OBUF2 REGF\[30\].RFW.BIT\[31\].FF/Q REGF\[30\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[31] sky130_fd_sc_hd__ebufn_2
XREGF\[9\].RFW.BIT\[19\].OBUF2 REGF\[9\].RFW.BIT\[19\].FF/Q REGF\[9\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[19] sky130_fd_sc_hd__ebufn_2
XREGF\[11\].RFW.BIT\[2\].OBUF1 REGF\[11\].RFW.BIT\[2\].FF/Q REGF\[11\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[2] sky130_fd_sc_hd__ebufn_2
Xfill_15_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_15_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_15_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XREGF\[14\].RFW.BIT\[27\].OBUF1 REGF\[14\].RFW.BIT\[27\].FF/Q REGF\[14\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[27] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[14\].OBUF2 REGF\[27\].RFW.BIT\[14\].FF/Q REGF\[27\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[14] sky130_fd_sc_hd__ebufn_2
Xfill_31_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_31_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[6\].RFW.BIT\[7\].OBUF2 REGF\[6\].RFW.BIT\[7\].FF/Q REGF\[6\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[7] sky130_fd_sc_hd__ebufn_2
XREGF\[1\].RFW.BIT\[17\].FF REGF\[1\].RFW.CG\[2\]/GCLK DW[17] VGND VGND VPWR VPWR
+ REGF\[1\].RFW.BIT\[17\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[1\].RFW.BIT\[1\].OBUF1 REGF\[1\].RFW.BIT\[1\].FF/Q REGF\[1\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[1] sky130_fd_sc_hd__ebufn_2
Xfill_61_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[7\].RFW.BIT\[11\].FF REGF\[7\].RFW.CG\[1\]/GCLK DW[11] VGND VGND VPWR VPWR
+ REGF\[7\].RFW.BIT\[11\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_54_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_47_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_3_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_3_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_3_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[17\].RFW.BIT\[12\].OBUF1 REGF\[17\].RFW.BIT\[12\].FF/Q REGF\[17\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[12] sky130_fd_sc_hd__ebufn_2
Xfill_2_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[18\].RFW.BIT\[28\].OBUF2 REGF\[18\].RFW.BIT\[28\].FF/Q REGF\[18\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[28] sky130_fd_sc_hd__ebufn_2
XREGF\[13\].RFW.BIT\[2\].OBUF1 REGF\[13\].RFW.BIT\[2\].FF/Q REGF\[13\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[2] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.BIT\[8\].OBUF2 REGF\[18\].RFW.BIT\[8\].FF/Q REGF\[18\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[8] sky130_fd_sc_hd__ebufn_2
Xtap_12_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[23\].RFW.BIT\[17\].OBUF2 REGF\[23\].RFW.BIT\[17\].FF/Q REGF\[23\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[17] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[30\].OBUF2 REGF\[24\].RFW.BIT\[30\].FF/Q REGF\[24\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[30] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[11\].FF REGF\[24\].RFW.CG\[1\]/GCLK DW[11] VGND VGND VPWR VPWR
+ REGF\[24\].RFW.BIT\[11\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_36_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_36_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[9\].RFW.BIT\[20\].OBUF2 REGF\[9\].RFW.BIT\[20\].FF/Q REGF\[9\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[20] sky130_fd_sc_hd__ebufn_2
Xfill_36_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[8\].RFW.BIT\[7\].OBUF2 REGF\[8\].RFW.BIT\[7\].FF/Q REGF\[8\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[7] sky130_fd_sc_hd__ebufn_2
Xfill_52_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[1\].RFW.BIT\[22\].OBUF1 REGF\[1\].RFW.BIT\[22\].FF/Q REGF\[1\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[22] sky130_fd_sc_hd__ebufn_2
Xfill_52_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_52_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.BIT\[1\].OBUF1 REGF\[3\].RFW.BIT\[1\].FF/Q REGF\[3\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[1] sky130_fd_sc_hd__ebufn_2
XREGF\[13\].RFW.BIT\[15\].OBUF1 REGF\[13\].RFW.BIT\[15\].FF/Q REGF\[13\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[15] sky130_fd_sc_hd__ebufn_2
XREGF\[11\].RFW.BIT\[6\].OBUF2 REGF\[11\].RFW.BIT\[6\].FF/Q REGF\[11\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[6] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.CGAND DEC2.D3.AND4/X WE VGND VGND VPWR VPWR REGF\[28\].RFW.CGAND/X
+ sky130_fd_sc_hd__and2_1
XREGF\[13\].RFW.BIT\[24\].FF REGF\[13\].RFW.CG\[3\]/GCLK DW[24] VGND VGND VPWR VPWR
+ REGF\[13\].RFW.BIT\[24\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_31_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[1\].RFW.BIT\[5\].OBUF2 REGF\[1\].RFW.BIT\[5\].FF/Q REGF\[1\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[5] sky130_fd_sc_hd__ebufn_2
Xfill_19_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[5\].RFW.BIT\[23\].OBUF2 REGF\[5\].RFW.BIT\[23\].FF/Q REGF\[5\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[23] sky130_fd_sc_hd__ebufn_2
XREGF\[15\].RFW.BIT\[2\].OBUF1 REGF\[15\].RFW.BIT\[2\].FF/Q REGF\[15\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[2] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.BIT\[16\].OBUF2 REGF\[17\].RFW.BIT\[16\].FF/Q REGF\[17\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[16] sky130_fd_sc_hd__ebufn_2
XREGF\[10\].RFW.BIT\[31\].OBUF1 REGF\[10\].RFW.BIT\[31\].FF/Q REGF\[10\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[31] sky130_fd_sc_hd__ebufn_2
Xfill_52_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_45_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[5\].RFW.BIT\[1\].OBUF1 REGF\[5\].RFW.BIT\[1\].FF/Q REGF\[5\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[1] sky130_fd_sc_hd__ebufn_2
XREGF\[14\].RFW.INV1\[0\] DEC0.D1.AND6/X VGND VGND VPWR VPWR REGF\[14\].RFW.INV1\[0\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_38_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[13\].RFW.BIT\[6\].OBUF2 REGF\[13\].RFW.BIT\[6\].FF/Q REGF\[13\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[6] sky130_fd_sc_hd__ebufn_2
XDEC2.D1.AND2 DEC2.D1.AND7/C DEC2.D1.AND7/A DEC2.D1.AND7/B DEC2.D1.AND7/D VGND VGND
+ VPWR VPWR DEC2.D1.AND2/X sky130_fd_sc_hd__and4bb_2
Xfill_22_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[8\].RFW.BIT\[17\].FF REGF\[8\].RFW.CG\[2\]/GCLK DW[17] VGND VGND VPWR VPWR
+ REGF\[8\].RFW.BIT\[17\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[1\].RFW.BIT\[26\].OBUF2 REGF\[1\].RFW.BIT\[26\].FF/Q REGF\[1\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[26] sky130_fd_sc_hd__ebufn_2
Xtap_10_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.BIT\[5\].OBUF2 REGF\[3\].RFW.BIT\[5\].FF/Q REGF\[3\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[5] sky130_fd_sc_hd__ebufn_2
XREGF\[13\].RFW.BIT\[19\].OBUF2 REGF\[13\].RFW.BIT\[19\].FF/Q REGF\[13\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[19] sky130_fd_sc_hd__ebufn_2
Xfill_47_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_47_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_47_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_47_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_3_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[17\].RFW.BIT\[2\].OBUF1 REGF\[17\].RFW.BIT\[2\].FF/Q REGF\[17\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[2] sky130_fd_sc_hd__ebufn_2
Xgenblk1.RFW0.BIT\[6\].OBUF1 genblk1.RFW0.TIE\[0\]/LO genblk1.RFW0.INV1\[0\]/Y VGND
+ VGND VPWR VPWR DA[6] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.BIT\[11\].OBUF2 REGF\[4\].RFW.BIT\[11\].FF/Q REGF\[4\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[11] sky130_fd_sc_hd__ebufn_2
Xfill_12_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[29\].RFW.BIT\[29\].OBUF1 REGF\[29\].RFW.BIT\[29\].FF/Q REGF\[29\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[29] sky130_fd_sc_hd__ebufn_2
XREGF\[7\].RFW.BIT\[1\].OBUF1 REGF\[7\].RFW.BIT\[1\].FF/Q REGF\[7\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[1] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.BIT\[2\].FF REGF\[19\].RFW.CG\[0\]/GCLK DW[2] VGND VGND VPWR VPWR
+ REGF\[19\].RFW.BIT\[2\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[25\].RFW.BIT\[17\].FF REGF\[25\].RFW.CG\[2\]/GCLK DW[17] VGND VGND VPWR VPWR
+ REGF\[25\].RFW.BIT\[17\].FF/Q sky130_fd_sc_hd__dfxtp_1
XDEC1.D2.AND4 DEC1.D2.AND7/A DEC1.D2.AND7/B DEC1.D2.AND7/C DEC1.D2.AND7/D VGND VGND
+ VPWR VPWR DEC1.D2.AND4/X sky130_fd_sc_hd__and4bb_2
XREGF\[10\].RFW.BIT\[0\].OBUF1 REGF\[10\].RFW.BIT\[0\].FF/Q REGF\[10\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[0] sky130_fd_sc_hd__ebufn_2
XREGF\[15\].RFW.BIT\[6\].OBUF2 REGF\[15\].RFW.BIT\[6\].FF/Q REGF\[15\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[6] sky130_fd_sc_hd__ebufn_2
Xfill_31_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_37_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_24_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_17_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.BIT\[4\].FF REGF\[18\].RFW.CG\[0\]/GCLK DW[4] VGND VGND VPWR VPWR
+ REGF\[18\].RFW.BIT\[4\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[5\].RFW.BIT\[5\].OBUF2 REGF\[5\].RFW.BIT\[5\].FF/Q REGF\[5\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[5] sky130_fd_sc_hd__ebufn_2
Xfill_9_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_9_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_9_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[19\].RFW.BIT\[2\].OBUF1 REGF\[19\].RFW.BIT\[2\].FF/Q REGF\[19\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[2] sky130_fd_sc_hd__ebufn_2
Xfill_50_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[13\].RFW.BIT\[20\].OBUF2 REGF\[13\].RFW.BIT\[20\].FF/Q REGF\[13\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[20] sky130_fd_sc_hd__ebufn_2
Xfill_17_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[17\].RFW.BIT\[6\].FF REGF\[17\].RFW.CG\[0\]/GCLK DW[6] VGND VGND VPWR VPWR
+ REGF\[17\].RFW.BIT\[6\].FF/Q sky130_fd_sc_hd__dfxtp_1
XDEC0.D3.ENBUF DEC0.D.AND3/X VGND VGND VPWR VPWR DEC0.D3.AND7/D sky130_fd_sc_hd__clkbuf_2
Xfill_33_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_33_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[24\].RFW.INV2\[2\] DEC1.D3.AND0/Y VGND VGND VPWR VPWR REGF\[24\].RFW.INV2\[2\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[9\].RFW.BIT\[1\].OBUF1 REGF\[9\].RFW.BIT\[1\].FF/Q REGF\[9\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[1] sky130_fd_sc_hd__ebufn_2
Xtap_10_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_58_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC0.D3.AND6 DEC0.D3.AND7/A DEC0.D3.AND7/B DEC0.D3.AND7/C DEC0.D3.AND7/D VGND VGND
+ VPWR VPWR DEC0.D3.AND6/X sky130_fd_sc_hd__and4b_2
XREGF\[28\].RFW.BIT\[17\].OBUF1 REGF\[28\].RFW.BIT\[17\].FF/Q REGF\[28\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[17] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.BIT\[30\].OBUF1 REGF\[29\].RFW.BIT\[30\].FF/Q REGF\[29\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[30] sky130_fd_sc_hd__ebufn_2
XREGF\[12\].RFW.BIT\[0\].OBUF1 REGF\[12\].RFW.BIT\[0\].FF/Q REGF\[12\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[0] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.BIT\[6\].OBUF2 REGF\[17\].RFW.BIT\[6\].FF/Q REGF\[17\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[6] sky130_fd_sc_hd__ebufn_2
Xfill_58_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_58_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_58_15 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[16\].RFW.BIT\[8\].FF REGF\[16\].RFW.CG\[1\]/GCLK DW[8] VGND VGND VPWR VPWR
+ REGF\[16\].RFW.BIT\[8\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_1_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[7\].RFW.BIT\[5\].OBUF2 REGF\[7\].RFW.BIT\[5\].FF/Q REGF\[7\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[5] sky130_fd_sc_hd__ebufn_2
Xfill_23_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.CG\[3\] CLK REGF\[3\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[3\].RFW.CG\[3\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_23_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[10\].RFW.BIT\[4\].OBUF2 REGF\[10\].RFW.BIT\[4\].FF/Q REGF\[10\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[4] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[25\].FF REGF\[5\].RFW.CG\[3\]/GCLK DW[25] VGND VGND VPWR VPWR
+ REGF\[5\].RFW.BIT\[25\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[11\].RFW.BIT\[15\].FF REGF\[11\].RFW.CG\[1\]/GCLK DW[15] VGND VGND VPWR VPWR
+ REGF\[11\].RFW.BIT\[15\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_22_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[20\].RFW.INV1\[3\] DEC0.D2.AND4/X VGND VGND VPWR VPWR REGF\[20\].RFW.INV1\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[30\].RFW.BIT\[22\].OBUF1 REGF\[30\].RFW.BIT\[22\].FF/Q REGF\[30\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[22] sky130_fd_sc_hd__ebufn_2
Xfill_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[29\].RFW.CG\[2\] CLK REGF\[29\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[29\].RFW.CG\[2\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[19\].RFW.BIT\[6\].OBUF2 REGF\[19\].RFW.BIT\[6\].FF/Q REGF\[19\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[6] sky130_fd_sc_hd__ebufn_2
XREGF\[14\].RFW.BIT\[0\].OBUF1 REGF\[14\].RFW.BIT\[0\].FF/Q REGF\[14\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[0] sky130_fd_sc_hd__ebufn_2
XREGF\[2\].RFW.CG\[0\] CLK REGF\[2\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[2\].RFW.CG\[0\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[21\].RFW.BIT\[9\].OBUF1 REGF\[21\].RFW.BIT\[9\].FF/Q REGF\[21\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[9] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.BIT\[8\].FF REGF\[29\].RFW.CG\[1\]/GCLK DW[8] VGND VGND VPWR VPWR
+ REGF\[29\].RFW.BIT\[8\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[9\].RFW.BIT\[5\].OBUF2 REGF\[9\].RFW.BIT\[5\].FF/Q REGF\[9\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[5] sky130_fd_sc_hd__ebufn_2
XREGF\[22\].RFW.BIT\[25\].FF REGF\[22\].RFW.CG\[3\]/GCLK DW[25] VGND VGND VPWR VPWR
+ REGF\[22\].RFW.BIT\[25\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_28_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[19\].RFW.INV2\[3\] DEC1.D2.AND3/X VGND VGND VPWR VPWR REGF\[19\].RFW.INV2\[3\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_44_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.BIT\[4\].OBUF2 REGF\[12\].RFW.BIT\[4\].FF/Q REGF\[12\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[4] sky130_fd_sc_hd__ebufn_2
Xfill_44_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_44_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_60_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_60_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_60_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_56_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.BIT\[26\].OBUF1 REGF\[6\].RFW.BIT\[26\].FF/Q REGF\[6\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[26] sky130_fd_sc_hd__ebufn_2
Xtap_49_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.BIT\[19\].OBUF1 REGF\[18\].RFW.BIT\[19\].FF/Q REGF\[18\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[19] sky130_fd_sc_hd__ebufn_2
XREGF\[2\].RFW.BIT\[3\].OBUF2 REGF\[2\].RFW.BIT\[3\].FF/Q REGF\[2\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[3] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[21\].OBUF1 REGF\[24\].RFW.BIT\[21\].FF/Q REGF\[24\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[21] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[0\].OBUF1 REGF\[16\].RFW.BIT\[0\].FF/Q REGF\[16\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[0] sky130_fd_sc_hd__ebufn_2
XREGF\[2\].RFW.BIT\[10\].FF REGF\[2\].RFW.CG\[1\]/GCLK DW[10] VGND VGND VPWR VPWR
+ REGF\[2\].RFW.BIT\[10\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[9\].RFW.BIT\[11\].OBUF1 REGF\[9\].RFW.BIT\[11\].FF/Q REGF\[9\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[11] sky130_fd_sc_hd__ebufn_2
XREGF\[23\].RFW.BIT\[9\].OBUF1 REGF\[23\].RFW.BIT\[9\].FF/Q REGF\[23\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[9] sky130_fd_sc_hd__ebufn_2
XREGF\[30\].RFW.BIT\[26\].OBUF2 REGF\[30\].RFW.BIT\[26\].FF/Q REGF\[30\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[26] sky130_fd_sc_hd__ebufn_2
Xfill_6_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_6_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[17\].RFW.CG\[2\] CLK REGF\[17\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[17\].RFW.CG\[2\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[14\].RFW.BIT\[4\].OBUF2 REGF\[14\].RFW.BIT\[4\].FF/Q REGF\[14\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[4] sky130_fd_sc_hd__ebufn_2
XREGF\[2\].RFW.BIT\[29\].OBUF1 REGF\[2\].RFW.BIT\[29\].FF/Q REGF\[2\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[29] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.BIT\[22\].OBUF2 REGF\[28\].RFW.BIT\[22\].FF/Q REGF\[28\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[22] sky130_fd_sc_hd__ebufn_2
Xfill_20_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_13_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[24\].OBUF1 REGF\[20\].RFW.BIT\[24\].FF/Q REGF\[20\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[24] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.BIT\[3\].OBUF2 REGF\[4\].RFW.BIT\[3\].FF/Q REGF\[4\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[3] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[14\].OBUF1 REGF\[5\].RFW.BIT\[14\].FF/Q REGF\[5\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[14] sky130_fd_sc_hd__ebufn_2
Xfill_30_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.BIT\[20\].OBUF1 REGF\[18\].RFW.BIT\[20\].FF/Q REGF\[18\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[20] sky130_fd_sc_hd__ebufn_2
Xtap_42_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.BIT\[0\].OBUF1 REGF\[18\].RFW.BIT\[0\].FF/Q REGF\[18\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[0] sky130_fd_sc_hd__ebufn_2
Xtap_28_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xtap_16_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_55_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_55_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.BIT\[15\].FF REGF\[18\].RFW.CG\[1\]/GCLK DW[15] VGND VGND VPWR VPWR
+ REGF\[18\].RFW.BIT\[15\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[25\].RFW.BIT\[9\].OBUF1 REGF\[25\].RFW.BIT\[9\].FF/Q REGF\[25\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[9] sky130_fd_sc_hd__ebufn_2
Xfill_55_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_55_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[30\].RFW.BIT\[20\].FF REGF\[30\].RFW.CG\[2\]/GCLK DW[20] VGND VGND VPWR VPWR
+ REGF\[30\].RFW.BIT\[20\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[24\].RFW.BIT\[25\].OBUF2 REGF\[24\].RFW.BIT\[25\].FF/Q REGF\[24\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[25] sky130_fd_sc_hd__ebufn_2
Xtap_61_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[16\].RFW.BIT\[4\].OBUF2 REGF\[16\].RFW.BIT\[4\].FF/Q REGF\[16\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[4] sky130_fd_sc_hd__ebufn_2
XREGF\[9\].RFW.BIT\[15\].OBUF2 REGF\[9\].RFW.BIT\[15\].FF/Q REGF\[9\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[15] sky130_fd_sc_hd__ebufn_2
Xfill_20_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[1\].RFW.BIT\[17\].OBUF1 REGF\[1\].RFW.BIT\[17\].FF/Q REGF\[1\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[17] sky130_fd_sc_hd__ebufn_2
XREGF\[2\].RFW.BIT\[30\].OBUF1 REGF\[2\].RFW.BIT\[30\].FF/Q REGF\[2\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[30] sky130_fd_sc_hd__ebufn_2
XREGF\[14\].RFW.BIT\[23\].OBUF1 REGF\[14\].RFW.BIT\[23\].FF/Q REGF\[14\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[23] sky130_fd_sc_hd__ebufn_2
Xfill_29_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_29_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[27\].RFW.BIT\[10\].OBUF2 REGF\[27\].RFW.BIT\[10\].FF/Q REGF\[27\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[10] sky130_fd_sc_hd__ebufn_2
Xfill_49_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[29\].RFW.BIT\[25\].FF REGF\[29\].RFW.CG\[3\]/GCLK DW[25] VGND VGND VPWR VPWR
+ REGF\[29\].RFW.BIT\[25\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[6\].RFW.BIT\[3\].OBUF2 REGF\[6\].RFW.BIT\[3\].FF/Q REGF\[6\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[3] sky130_fd_sc_hd__ebufn_2
XREGF\[6\].RFW.INV2\[1\] DEC1.D0.AND6/X VGND VGND VPWR VPWR REGF\[6\].RFW.INV2\[1\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_4_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_45_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[28\].OBUF2 REGF\[20\].RFW.BIT\[28\].FF/Q REGF\[20\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[28] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[9\].OBUF1 REGF\[27\].RFW.BIT\[9\].FF/Q REGF\[27\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[9] sky130_fd_sc_hd__ebufn_2
XREGF\[6\].RFW.BIT\[31\].OBUF2 REGF\[6\].RFW.BIT\[31\].FF/Q REGF\[6\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[31] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[18\].OBUF2 REGF\[5\].RFW.BIT\[18\].FF/Q REGF\[5\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[18] sky130_fd_sc_hd__ebufn_2
XREGF\[3\].RFW.BIT\[16\].FF REGF\[3\].RFW.CG\[2\]/GCLK DW[16] VGND VGND VPWR VPWR
+ REGF\[3\].RFW.BIT\[16\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[18\].RFW.BIT\[24\].OBUF2 REGF\[18\].RFW.BIT\[24\].FF/Q REGF\[18\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[24] sky130_fd_sc_hd__ebufn_2
Xfill_25_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[9\].RFW.BIT\[10\].FF REGF\[9\].RFW.CG\[1\]/GCLK DW[10] VGND VGND VPWR VPWR
+ REGF\[9\].RFW.BIT\[10\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_8_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.BIT\[4\].OBUF2 REGF\[18\].RFW.BIT\[4\].FF/Q REGF\[18\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[4] sky130_fd_sc_hd__ebufn_2
XREGF\[10\].RFW.BIT\[26\].OBUF1 REGF\[10\].RFW.BIT\[26\].FF/Q REGF\[10\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[26] sky130_fd_sc_hd__ebufn_2
XREGF\[23\].RFW.BIT\[13\].OBUF2 REGF\[23\].RFW.BIT\[13\].FF/Q REGF\[23\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[13] sky130_fd_sc_hd__ebufn_2
Xfill_41_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_41_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[27\].RFW.CGAND DEC2.D3.AND3/X WE VGND VGND VPWR VPWR REGF\[27\].RFW.CGAND/X
+ sky130_fd_sc_hd__and2_1
XREGF\[20\].RFW.BIT\[7\].OBUF1 REGF\[20\].RFW.BIT\[7\].FF/Q REGF\[20\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[7] sky130_fd_sc_hd__ebufn_2
Xtap_40_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[8\].RFW.BIT\[3\].OBUF2 REGF\[8\].RFW.BIT\[3\].FF/Q REGF\[8\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[3] sky130_fd_sc_hd__ebufn_2
Xtap_26_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[13\].RFW.BIT\[11\].OBUF1 REGF\[13\].RFW.BIT\[11\].FF/Q REGF\[13\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[11] sky130_fd_sc_hd__ebufn_2
XREGF\[2\].RFW.INV1\[2\] DEC0.D0.AND2/X VGND VGND VPWR VPWR REGF\[2\].RFW.INV1\[2\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[20\].RFW.BIT\[16\].FF REGF\[20\].RFW.CG\[2\]/GCLK DW[16] VGND VGND VPWR VPWR
+ REGF\[20\].RFW.BIT\[16\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[11\].RFW.BIT\[2\].OBUF2 REGF\[11\].RFW.BIT\[2\].FF/Q REGF\[11\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[2] sky130_fd_sc_hd__ebufn_2
Xfill_15_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_15_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[26\].RFW.BIT\[10\].FF REGF\[26\].RFW.CG\[1\]/GCLK DW[10] VGND VGND VPWR VPWR
+ REGF\[26\].RFW.BIT\[10\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_15_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XREGF\[13\].RFW.BIT\[1\].FF REGF\[13\].RFW.CG\[0\]/GCLK DW[1] VGND VGND VPWR VPWR
+ REGF\[13\].RFW.BIT\[1\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[29\].RFW.BIT\[9\].OBUF1 REGF\[29\].RFW.BIT\[9\].FF/Q REGF\[29\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[9] sky130_fd_sc_hd__ebufn_2
XREGF\[14\].RFW.BIT\[27\].OBUF2 REGF\[14\].RFW.BIT\[27\].FF/Q REGF\[14\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[27] sky130_fd_sc_hd__ebufn_2
Xfill_31_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_31_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[1\].RFW.BIT\[1\].OBUF2 REGF\[1\].RFW.BIT\[1\].FF/Q REGF\[1\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[1] sky130_fd_sc_hd__ebufn_2
XREGF\[22\].RFW.INV1\[0\] DEC0.D2.AND6/X VGND VGND VPWR VPWR REGF\[22\].RFW.INV1\[0\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_61_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_54_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_47_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_3_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_3_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_3_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[15\].RFW.BIT\[23\].FF REGF\[15\].RFW.CG\[2\]/GCLK DW[23] VGND VGND VPWR VPWR
+ REGF\[15\].RFW.BIT\[23\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[17\].RFW.BIT\[12\].OBUF2 REGF\[17\].RFW.BIT\[12\].FF/Q REGF\[17\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[12] sky130_fd_sc_hd__ebufn_2
XREGF\[12\].RFW.BIT\[3\].FF REGF\[12\].RFW.CG\[0\]/GCLK DW[3] VGND VGND VPWR VPWR
+ REGF\[12\].RFW.BIT\[3\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[31\].RFW.BIT\[26\].FF REGF\[31\].RFW.CG\[3\]/GCLK DW[26] VGND VGND VPWR VPWR
+ REGF\[31\].RFW.BIT\[26\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_2_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[22\].RFW.BIT\[7\].OBUF1 REGF\[22\].RFW.BIT\[7\].FF/Q REGF\[22\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[7] sky130_fd_sc_hd__ebufn_2
XREGF\[13\].RFW.BIT\[2\].OBUF2 REGF\[13\].RFW.BIT\[2\].FF/Q REGF\[13\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[2] sky130_fd_sc_hd__ebufn_2
XREGF\[11\].RFW.BIT\[5\].FF REGF\[11\].RFW.CG\[0\]/GCLK DW[5] VGND VGND VPWR VPWR
+ REGF\[11\].RFW.BIT\[5\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_12_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_36_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_52_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_52_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_52_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[1\].RFW.BIT\[22\].OBUF2 REGF\[1\].RFW.BIT\[22\].FF/Q REGF\[1\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[22] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[1\].FF REGF\[26\].RFW.CG\[0\]/GCLK DW[1] VGND VGND VPWR VPWR
+ REGF\[26\].RFW.BIT\[1\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[3\].RFW.BIT\[1\].OBUF2 REGF\[3\].RFW.BIT\[1\].FF/Q REGF\[3\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[1] sky130_fd_sc_hd__ebufn_2
XREGF\[13\].RFW.BIT\[15\].OBUF2 REGF\[13\].RFW.BIT\[15\].FF/Q REGF\[13\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[15] sky130_fd_sc_hd__ebufn_2
XREGF\[10\].RFW.BIT\[7\].FF REGF\[10\].RFW.CG\[0\]/GCLK DW[7] VGND VGND VPWR VPWR
+ REGF\[10\].RFW.BIT\[7\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_31_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.BIT\[29\].OBUF1 REGF\[31\].RFW.BIT\[29\].FF/Q REGF\[31\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[29] sky130_fd_sc_hd__ebufn_2
Xtap_24_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgenblk1.RFW0.BIT\[2\].OBUF1 genblk1.RFW0.TIE\[0\]/LO genblk1.RFW0.INV1\[0\]/Y VGND
+ VGND VPWR VPWR DA[2] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[7\].OBUF1 REGF\[24\].RFW.BIT\[7\].FF/Q REGF\[24\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[7] sky130_fd_sc_hd__ebufn_2
XREGF\[25\].RFW.BIT\[3\].FF REGF\[25\].RFW.CG\[0\]/GCLK DW[3] VGND VGND VPWR VPWR
+ REGF\[25\].RFW.BIT\[3\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[29\].RFW.BIT\[25\].OBUF1 REGF\[29\].RFW.BIT\[25\].FF/Q REGF\[29\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[25] sky130_fd_sc_hd__ebufn_2
XREGF\[15\].RFW.BIT\[2\].OBUF2 REGF\[15\].RFW.BIT\[2\].FF/Q REGF\[15\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[2] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.INV1\[1\] DEC0.D2.AND1/X VGND VGND VPWR VPWR REGF\[17\].RFW.INV1\[1\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[24\].RFW.BIT\[5\].FF REGF\[24\].RFW.CG\[0\]/GCLK DW[5] VGND VGND VPWR VPWR
+ REGF\[24\].RFW.BIT\[5\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[10\].RFW.BIT\[31\].OBUF2 REGF\[10\].RFW.BIT\[31\].FF/Q REGF\[10\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[31] sky130_fd_sc_hd__ebufn_2
Xfill_52_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_45_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[5\].RFW.BIT\[1\].OBUF2 REGF\[5\].RFW.BIT\[1\].FF/Q REGF\[5\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[1] sky130_fd_sc_hd__ebufn_2
Xfill_38_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[27\].RFW.BIT\[16\].FF REGF\[27\].RFW.CG\[2\]/GCLK DW[16] VGND VGND VPWR VPWR
+ REGF\[27\].RFW.BIT\[16\].FF/Q sky130_fd_sc_hd__dfxtp_1
XDEC2.D1.AND3 DEC2.D1.AND7/C DEC2.D1.AND7/B DEC2.D1.AND7/A DEC2.D1.AND7/D VGND VGND
+ VPWR VPWR DEC2.D1.AND3/X sky130_fd_sc_hd__and4b_2
XREGF\[23\].RFW.BIT\[7\].FF REGF\[23\].RFW.CG\[0\]/GCLK DW[7] VGND VGND VPWR VPWR
+ REGF\[23\].RFW.BIT\[7\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[25\].RFW.BIT\[28\].OBUF1 REGF\[25\].RFW.BIT\[28\].FF/Q REGF\[25\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[28] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[7\].OBUF1 REGF\[26\].RFW.BIT\[7\].FF/Q REGF\[26\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[7] sky130_fd_sc_hd__ebufn_2
XREGF\[30\].RFW.BIT\[17\].OBUF1 REGF\[30\].RFW.BIT\[17\].FF/Q REGF\[30\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[17] sky130_fd_sc_hd__ebufn_2
XREGF\[31\].RFW.BIT\[30\].OBUF1 REGF\[31\].RFW.BIT\[30\].FF/Q REGF\[31\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[30] sky130_fd_sc_hd__ebufn_2
Xtap_10_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[9\].RFW.BIT\[2\].FF REGF\[9\].RFW.CG\[0\]/GCLK DW[2] VGND VGND VPWR VPWR REGF\[9\].RFW.BIT\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xfill_47_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_47_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[16\].RFW.BIT\[29\].FF REGF\[16\].RFW.CG\[3\]/GCLK DW[29] VGND VGND VPWR VPWR
+ REGF\[16\].RFW.BIT\[29\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_47_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XREGF\[12\].RFW.BIT\[31\].FF REGF\[12\].RFW.CG\[3\]/GCLK DW[31] VGND VGND VPWR VPWR
+ REGF\[12\].RFW.BIT\[31\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_3_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[22\].RFW.BIT\[9\].FF REGF\[22\].RFW.CG\[1\]/GCLK DW[9] VGND VGND VPWR VPWR
+ REGF\[22\].RFW.BIT\[9\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[28\].RFW.BIT\[13\].OBUF1 REGF\[28\].RFW.BIT\[13\].FF/Q REGF\[28\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[13] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.BIT\[2\].OBUF2 REGF\[17\].RFW.BIT\[2\].FF/Q REGF\[17\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[2] sky130_fd_sc_hd__ebufn_2
Xgenblk1.RFW0.BIT\[6\].OBUF2 genblk1.RFW0.TIE\[4\]/LO genblk1.RFW0.INV2\[0\]/Y VGND
+ VGND VPWR VPWR DB[6] sky130_fd_sc_hd__ebufn_2
Xfill_12_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_12_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[8\].RFW.BIT\[4\].FF REGF\[8\].RFW.CG\[0\]/GCLK DW[4] VGND VGND VPWR VPWR REGF\[8\].RFW.BIT\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[29\].RFW.BIT\[29\].OBUF2 REGF\[29\].RFW.BIT\[29\].FF/Q REGF\[29\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[29] sky130_fd_sc_hd__ebufn_2
XREGF\[7\].RFW.BIT\[1\].OBUF2 REGF\[7\].RFW.BIT\[1\].FF/Q REGF\[7\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[1] sky130_fd_sc_hd__ebufn_2
XDEC1.D2.AND5 DEC1.D2.AND7/B DEC1.D2.AND7/A DEC1.D2.AND7/C DEC1.D2.AND7/D VGND VGND
+ VPWR VPWR DEC1.D2.AND5/X sky130_fd_sc_hd__and4b_2
XREGF\[10\].RFW.BIT\[0\].OBUF2 REGF\[10\].RFW.BIT\[0\].FF/Q REGF\[10\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[0] sky130_fd_sc_hd__ebufn_2
Xfill_31_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[25\].RFW.CG\[1\] CLK REGF\[25\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[25\].RFW.CG\[1\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_37_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_37_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_24_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_17_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[19\].RFW.BIT\[27\].OBUF1 REGF\[19\].RFW.BIT\[27\].FF/Q REGF\[19\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[27] sky130_fd_sc_hd__ebufn_2
XREGF\[7\].RFW.BIT\[6\].FF REGF\[7\].RFW.CG\[0\]/GCLK DW[6] VGND VGND VPWR VPWR REGF\[7\].RFW.BIT\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xfill_0_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_53_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[28\].RFW.BIT\[7\].OBUF1 REGF\[28\].RFW.BIT\[7\].FF/Q REGF\[28\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[7] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[16\].OBUF1 REGF\[24\].RFW.BIT\[16\].FF/Q REGF\[24\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[16] sky130_fd_sc_hd__ebufn_2
Xfill_9_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_9_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_9_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[11\].RFW.INV2\[2\] DEC1.D1.AND3/X VGND VGND VPWR VPWR REGF\[11\].RFW.INV2\[2\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XREGF\[27\].RFW.INV2\[3\] DEC1.D3.AND3/X VGND VGND VPWR VPWR REGF\[27\].RFW.INV2\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[19\].RFW.BIT\[2\].OBUF2 REGF\[19\].RFW.BIT\[2\].FF/Q REGF\[19\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[2] sky130_fd_sc_hd__ebufn_2
Xfill_50_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[6\].RFW.BIT\[8\].FF REGF\[6\].RFW.CG\[1\]/GCLK DW[8] VGND VGND VPWR VPWR REGF\[6\].RFW.BIT\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xfill_43_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[7\].RFW.BIT\[24\].FF REGF\[7\].RFW.CG\[3\]/GCLK DW[24] VGND VGND VPWR VPWR
+ REGF\[7\].RFW.BIT\[24\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[21\].RFW.BIT\[5\].OBUF1 REGF\[21\].RFW.BIT\[5\].FF/Q REGF\[21\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[5] sky130_fd_sc_hd__ebufn_2
XREGF\[13\].RFW.BIT\[14\].FF REGF\[13\].RFW.CG\[1\]/GCLK DW[14] VGND VGND VPWR VPWR
+ REGF\[13\].RFW.BIT\[14\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_33_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[9\].RFW.BIT\[1\].OBUF2 REGF\[9\].RFW.BIT\[1\].FF/Q REGF\[9\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[1] sky130_fd_sc_hd__ebufn_2
Xtap_10_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_58_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC0.D3.AND7 DEC0.D3.AND7/A DEC0.D3.AND7/B DEC0.D3.AND7/C DEC0.D3.AND7/D VGND VGND
+ VPWR VPWR DEC0.D3.AND7/X sky130_fd_sc_hd__and4_2
XREGF\[28\].RFW.BIT\[17\].OBUF2 REGF\[28\].RFW.BIT\[17\].FF/Q REGF\[28\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[17] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.BIT\[30\].OBUF2 REGF\[29\].RFW.BIT\[30\].FF/Q REGF\[29\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[30] sky130_fd_sc_hd__ebufn_2
XREGF\[12\].RFW.BIT\[0\].OBUF2 REGF\[12\].RFW.BIT\[0\].FF/Q REGF\[12\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[0] sky130_fd_sc_hd__ebufn_2
XREGF\[20\].RFW.BIT\[19\].OBUF1 REGF\[20\].RFW.BIT\[19\].FF/Q REGF\[20\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[19] sky130_fd_sc_hd__ebufn_2
Xfill_58_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_58_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_58_16 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.BIT\[22\].OBUF1 REGF\[6\].RFW.BIT\[22\].FF/Q REGF\[6\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[22] sky130_fd_sc_hd__ebufn_2
Xtap_1_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.BIT\[15\].OBUF1 REGF\[18\].RFW.BIT\[15\].FF/Q REGF\[18\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[15] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[24\].FF REGF\[24\].RFW.CG\[3\]/GCLK DW[24] VGND VGND VPWR VPWR
+ REGF\[24\].RFW.BIT\[24\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_23_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_23_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_23_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[13\].RFW.CG\[1\] CLK REGF\[13\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[13\].RFW.CG\[1\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[23\].RFW.BIT\[5\].OBUF1 REGF\[23\].RFW.BIT\[5\].FF/Q REGF\[23\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[5] sky130_fd_sc_hd__ebufn_2
Xfill_22_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[30\].RFW.BIT\[22\].OBUF2 REGF\[30\].RFW.BIT\[22\].FF/Q REGF\[30\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[22] sky130_fd_sc_hd__ebufn_2
Xfill_15_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[19\].RFW.BIT\[31\].FF REGF\[19\].RFW.CG\[3\]/GCLK DW[31] VGND VGND VPWR VPWR
+ REGF\[19\].RFW.BIT\[31\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[14\].RFW.BIT\[0\].OBUF2 REGF\[14\].RFW.BIT\[0\].FF/Q REGF\[14\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[0] sky130_fd_sc_hd__ebufn_2
XREGF\[2\].RFW.BIT\[25\].OBUF1 REGF\[2\].RFW.BIT\[25\].FF/Q REGF\[2\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[25] sky130_fd_sc_hd__ebufn_2
XREGF\[14\].RFW.BIT\[18\].OBUF1 REGF\[14\].RFW.BIT\[18\].FF/Q REGF\[14\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[18] sky130_fd_sc_hd__ebufn_2
XREGF\[15\].RFW.BIT\[31\].OBUF1 REGF\[15\].RFW.BIT\[31\].FF/Q REGF\[15\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[31] sky130_fd_sc_hd__ebufn_2
XREGF\[20\].RFW.BIT\[20\].OBUF1 REGF\[20\].RFW.BIT\[20\].FF/Q REGF\[20\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[20] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.BIT\[9\].OBUF2 REGF\[21\].RFW.BIT\[9\].FF/Q REGF\[21\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[9] sky130_fd_sc_hd__ebufn_2
Xfill_28_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[5\].RFW.BIT\[10\].OBUF1 REGF\[5\].RFW.BIT\[10\].FF/Q REGF\[5\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[10] sky130_fd_sc_hd__ebufn_2
Xfill_44_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDEC2.D2.ABUF\[2\] RW[2] VGND VGND VPWR VPWR DEC2.D2.AND7/C sky130_fd_sc_hd__clkbuf_2
Xfill_60_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_60_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_60_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_56_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.BIT\[26\].OBUF2 REGF\[6\].RFW.BIT\[26\].FF/Q REGF\[6\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[26] sky130_fd_sc_hd__ebufn_2
XREGF\[25\].RFW.BIT\[5\].OBUF1 REGF\[25\].RFW.BIT\[5\].FF/Q REGF\[25\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[5] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.BIT\[19\].OBUF2 REGF\[18\].RFW.BIT\[19\].FF/Q REGF\[18\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[19] sky130_fd_sc_hd__ebufn_2
Xtap_49_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[24\].RFW.BIT\[21\].OBUF2 REGF\[24\].RFW.BIT\[21\].FF/Q REGF\[24\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[21] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[0\].OBUF2 REGF\[16\].RFW.BIT\[0\].FF/Q REGF\[16\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[0] sky130_fd_sc_hd__ebufn_2
Xfill_18_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[9\].RFW.BIT\[11\].OBUF2 REGF\[9\].RFW.BIT\[11\].FF/Q REGF\[9\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[11] sky130_fd_sc_hd__ebufn_2
XREGF\[10\].RFW.BIT\[22\].FF REGF\[10\].RFW.CG\[2\]/GCLK DW[22] VGND VGND VPWR VPWR
+ REGF\[10\].RFW.BIT\[22\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_34_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[1\].RFW.BIT\[13\].OBUF1 REGF\[1\].RFW.BIT\[13\].FF/Q REGF\[1\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[13] sky130_fd_sc_hd__ebufn_2
XREGF\[23\].RFW.BIT\[9\].OBUF2 REGF\[23\].RFW.BIT\[9\].FF/Q REGF\[23\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[9] sky130_fd_sc_hd__ebufn_2
Xfill_6_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_6_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_6_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgenblk1.RFW0.TIE\[6\] VGND VGND VPWR VPWR genblk1.RFW0.TIE\[6\]/HI genblk1.RFW0.TIE\[6\]/LO
+ sky130_fd_sc_hd__conb_1
XDEC0.D2.ENBUF DEC0.D.AND2/X VGND VGND VPWR VPWR DEC0.D2.AND7/D sky130_fd_sc_hd__clkbuf_2
XREGF\[2\].RFW.BIT\[29\].OBUF2 REGF\[2\].RFW.BIT\[29\].FF/Q REGF\[2\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[29] sky130_fd_sc_hd__ebufn_2
Xfill_20_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfill_13_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[20\].RFW.BIT\[24\].OBUF2 REGF\[20\].RFW.BIT\[24\].FF/Q REGF\[20\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[24] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[5\].OBUF1 REGF\[27\].RFW.BIT\[5\].FF/Q REGF\[27\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[5] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[14\].OBUF2 REGF\[5\].RFW.BIT\[14\].FF/Q REGF\[5\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[14] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.CGAND DEC2.D3.AND2/X WE VGND VGND VPWR VPWR REGF\[26\].RFW.CGAND/X
+ sky130_fd_sc_hd__and2_1
XREGF\[18\].RFW.BIT\[20\].OBUF2 REGF\[18\].RFW.BIT\[20\].FF/Q REGF\[18\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[20] sky130_fd_sc_hd__ebufn_2
Xtap_42_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.BIT\[0\].OBUF2 REGF\[18\].RFW.BIT\[0\].FF/Q REGF\[18\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[0] sky130_fd_sc_hd__ebufn_2
Xtap_28_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[10\].RFW.BIT\[22\].OBUF1 REGF\[10\].RFW.BIT\[22\].FF/Q REGF\[10\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[22] sky130_fd_sc_hd__ebufn_2
Xfill_39_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_39_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xtap_16_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[0\].FF REGF\[20\].RFW.CG\[0\]/GCLK DW[0] VGND VGND VPWR VPWR
+ REGF\[20\].RFW.BIT\[0\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_55_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[25\].RFW.BIT\[9\].OBUF2 REGF\[25\].RFW.BIT\[9\].FF/Q REGF\[25\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[9] sky130_fd_sc_hd__ebufn_2
Xfill_55_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_55_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[3\].OBUF1 REGF\[20\].RFW.BIT\[3\].FF/Q REGF\[20\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[3] sky130_fd_sc_hd__ebufn_2
Xtap_32_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[5\].RFW.BIT\[15\].FF REGF\[5\].RFW.CG\[1\]/GCLK DW[15] VGND VGND VPWR VPWR
+ REGF\[5\].RFW.BIT\[15\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_61_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[30\].RFW.INV1\[0\] DEC0.D3.AND6/X VGND VGND VPWR VPWR REGF\[30\].RFW.INV1\[0\]/Y
+ sky130_fd_sc_hd__inv_4
Xtap_54_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[9\].RFW.INV2\[2\] DEC1.D1.AND1/X VGND VGND VPWR VPWR REGF\[9\].RFW.INV2\[2\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_20_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_20_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[1\].RFW.BIT\[17\].OBUF2 REGF\[1\].RFW.BIT\[17\].FF/Q REGF\[1\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[17] sky130_fd_sc_hd__ebufn_2
XREGF\[2\].RFW.BIT\[30\].OBUF2 REGF\[2\].RFW.BIT\[30\].FF/Q REGF\[2\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[30] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.BIT\[5\].OBUF1 REGF\[29\].RFW.BIT\[5\].FF/Q REGF\[29\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[5] sky130_fd_sc_hd__ebufn_2
XREGF\[14\].RFW.BIT\[23\].OBUF2 REGF\[14\].RFW.BIT\[23\].FF/Q REGF\[14\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[23] sky130_fd_sc_hd__ebufn_2
Xfill_29_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_29_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_45_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_45_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[29\].RFW.INV2\[0\] DEC1.D3.AND5/X VGND VGND VPWR VPWR REGF\[29\].RFW.INV2\[0\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_61_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[22\].RFW.BIT\[15\].FF REGF\[22\].RFW.CG\[1\]/GCLK DW[15] VGND VGND VPWR VPWR
+ REGF\[22\].RFW.BIT\[15\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[27\].RFW.BIT\[9\].OBUF2 REGF\[27\].RFW.BIT\[9\].FF/Q REGF\[27\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[9] sky130_fd_sc_hd__ebufn_2
XREGF\[22\].RFW.BIT\[3\].OBUF1 REGF\[22\].RFW.BIT\[3\].FF/Q REGF\[22\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[3] sky130_fd_sc_hd__ebufn_2
Xfill_9_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[11\].RFW.BIT\[28\].FF REGF\[11\].RFW.CG\[3\]/GCLK DW[28] VGND VGND VPWR VPWR
+ REGF\[11\].RFW.BIT\[28\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[10\].RFW.BIT\[26\].OBUF2 REGF\[10\].RFW.BIT\[26\].FF/Q REGF\[10\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[26] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.INV1\[3\] DEC0.D0.AND5/X VGND VGND VPWR VPWR REGF\[5\].RFW.INV1\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[17\].RFW.BIT\[22\].FF REGF\[17\].RFW.CG\[2\]/GCLK DW[22] VGND VGND VPWR VPWR
+ REGF\[17\].RFW.BIT\[22\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_41_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.BIT\[1\].FF REGF\[3\].RFW.CG\[0\]/GCLK DW[1] VGND VGND VPWR VPWR REGF\[3\].RFW.BIT\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[20\].RFW.BIT\[7\].OBUF2 REGF\[20\].RFW.BIT\[7\].FF/Q REGF\[20\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[7] sky130_fd_sc_hd__ebufn_2
Xtap_40_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_19_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[13\].RFW.BIT\[11\].OBUF2 REGF\[13\].RFW.BIT\[11\].FF/Q REGF\[13\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[11] sky130_fd_sc_hd__ebufn_2
XREGF\[25\].RFW.INV1\[1\] DEC0.D3.AND1/X VGND VGND VPWR VPWR REGF\[25\].RFW.INV1\[1\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[2\].RFW.BIT\[3\].FF REGF\[2\].RFW.CG\[0\]/GCLK DW[3] VGND VGND VPWR VPWR REGF\[2\].RFW.BIT\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XREGF\[31\].RFW.BIT\[4\].FF REGF\[31\].RFW.CG\[0\]/GCLK DW[4] VGND VGND VPWR VPWR
+ REGF\[31\].RFW.BIT\[4\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[31\].RFW.BIT\[25\].OBUF1 REGF\[31\].RFW.BIT\[25\].FF/Q REGF\[31\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[25] sky130_fd_sc_hd__ebufn_2
Xfill_15_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_15_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_15_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_15_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[29\].RFW.BIT\[9\].OBUF2 REGF\[29\].RFW.BIT\[9\].FF/Q REGF\[29\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[9] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[3\].OBUF1 REGF\[24\].RFW.BIT\[3\].FF/Q REGF\[24\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[3] sky130_fd_sc_hd__ebufn_2
Xfill_31_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_31_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_31_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_31_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XREGF\[29\].RFW.BIT\[21\].OBUF1 REGF\[29\].RFW.BIT\[21\].FF/Q REGF\[29\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[21] sky130_fd_sc_hd__ebufn_2
Xfill_61_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_54_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[30\].RFW.BIT\[6\].FF REGF\[30\].RFW.CG\[0\]/GCLK DW[6] VGND VGND VPWR VPWR
+ REGF\[30\].RFW.BIT\[6\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[1\].RFW.BIT\[5\].FF REGF\[1\].RFW.CG\[0\]/GCLK DW[5] VGND VGND VPWR VPWR REGF\[1\].RFW.BIT\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xfill_3_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_47_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_2_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[22\].RFW.BIT\[7\].OBUF2 REGF\[22\].RFW.BIT\[7\].FF/Q REGF\[22\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[7] sky130_fd_sc_hd__ebufn_2
XREGF\[2\].RFW.BIT\[23\].FF REGF\[2\].RFW.CG\[2\]/GCLK DW[23] VGND VGND VPWR VPWR
+ REGF\[2\].RFW.BIT\[23\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[7\].RFW.BIT\[29\].OBUF1 REGF\[7\].RFW.BIT\[29\].FF/Q REGF\[7\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[29] sky130_fd_sc_hd__ebufn_2
XREGF\[22\].RFW.CG\[3\] CLK REGF\[22\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[22\].RFW.CG\[3\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[30\].RFW.BIT\[10\].FF REGF\[30\].RFW.CG\[1\]/GCLK DW[10] VGND VGND VPWR VPWR
+ REGF\[30\].RFW.BIT\[10\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[25\].RFW.BIT\[24\].OBUF1 REGF\[25\].RFW.BIT\[24\].FF/Q REGF\[25\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[24] sky130_fd_sc_hd__ebufn_2
Xfill_36_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[30\].RFW.BIT\[13\].OBUF1 REGF\[30\].RFW.BIT\[13\].FF/Q REGF\[30\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[13] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[3\].OBUF1 REGF\[26\].RFW.BIT\[3\].FF/Q REGF\[26\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[3] sky130_fd_sc_hd__ebufn_2
Xfill_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_52_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[29\].RFW.BIT\[15\].FF REGF\[29\].RFW.CG\[1\]/GCLK DW[15] VGND VGND VPWR VPWR
+ REGF\[29\].RFW.BIT\[15\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_31_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.BIT\[29\].OBUF2 REGF\[31\].RFW.BIT\[29\].FF/Q REGF\[31\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[29] sky130_fd_sc_hd__ebufn_2
Xgenblk1.RFW0.BIT\[2\].OBUF2 genblk1.RFW0.TIE\[4\]/LO genblk1.RFW0.INV2\[0\]/Y VGND
+ VGND VPWR VPWR DB[2] sky130_fd_sc_hd__ebufn_2
Xtap_24_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[21\].RFW.CG\[0\] CLK REGF\[21\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[21\].RFW.CG\[0\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[24\].RFW.BIT\[7\].OBUF2 REGF\[24\].RFW.BIT\[7\].FF/Q REGF\[24\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[7] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.BIT\[25\].OBUF2 REGF\[29\].RFW.BIT\[25\].FF/Q REGF\[29\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[25] sky130_fd_sc_hd__ebufn_2
Xfill_26_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[21\].RFW.BIT\[27\].OBUF1 REGF\[21\].RFW.BIT\[27\].FF/Q REGF\[21\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[27] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.BIT\[28\].FF REGF\[18\].RFW.CG\[3\]/GCLK DW[28] VGND VGND VPWR VPWR
+ REGF\[18\].RFW.BIT\[28\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[14\].RFW.BIT\[30\].FF REGF\[14\].RFW.CG\[3\]/GCLK DW[30] VGND VGND VPWR VPWR
+ REGF\[14\].RFW.BIT\[30\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_42_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[7\].RFW.BIT\[30\].OBUF1 REGF\[7\].RFW.BIT\[30\].FF/Q REGF\[7\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[30] sky130_fd_sc_hd__ebufn_2
XREGF\[6\].RFW.BIT\[17\].OBUF1 REGF\[6\].RFW.BIT\[17\].FF/Q REGF\[6\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[17] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.BIT\[23\].OBUF1 REGF\[19\].RFW.BIT\[23\].FF/Q REGF\[19\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[23] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.BIT\[3\].OBUF1 REGF\[28\].RFW.BIT\[3\].FF/Q REGF\[28\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[3] sky130_fd_sc_hd__ebufn_2
Xfill_52_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[24\].RFW.BIT\[12\].OBUF1 REGF\[24\].RFW.BIT\[12\].FF/Q REGF\[24\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[12] sky130_fd_sc_hd__ebufn_2
Xfill_45_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_38_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[10\].RFW.CG\[3\] CLK REGF\[10\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[10\].RFW.CG\[3\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XDEC2.D1.AND4 DEC2.D1.AND7/A DEC2.D1.AND7/B DEC2.D1.AND7/C DEC2.D1.AND7/D VGND VGND
+ VPWR VPWR DEC2.D1.AND4/X sky130_fd_sc_hd__and4bb_2
XREGF\[25\].RFW.BIT\[28\].OBUF2 REGF\[25\].RFW.BIT\[28\].FF/Q REGF\[25\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[28] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[7\].OBUF2 REGF\[26\].RFW.BIT\[7\].FF/Q REGF\[26\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[7] sky130_fd_sc_hd__ebufn_2
XREGF\[30\].RFW.BIT\[17\].OBUF2 REGF\[30\].RFW.BIT\[17\].FF/Q REGF\[30\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[17] sky130_fd_sc_hd__ebufn_2
XREGF\[31\].RFW.BIT\[30\].OBUF2 REGF\[31\].RFW.BIT\[30\].FF/Q REGF\[31\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[30] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.BIT\[1\].OBUF1 REGF\[21\].RFW.BIT\[1\].FF/Q REGF\[21\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[1] sky130_fd_sc_hd__ebufn_2
Xtap_10_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_47_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_47_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[15\].RFW.BIT\[26\].OBUF1 REGF\[15\].RFW.BIT\[26\].FF/Q REGF\[15\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[26] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.BIT\[13\].OBUF2 REGF\[28\].RFW.BIT\[13\].FF/Q REGF\[28\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[13] sky130_fd_sc_hd__ebufn_2
Xtap_24_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[15\].OBUF1 REGF\[20\].RFW.BIT\[15\].FF/Q REGF\[20\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[15] sky130_fd_sc_hd__ebufn_2
Xtap_40_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[3\].RFW.BIT\[29\].FF REGF\[3\].RFW.CG\[3\]/GCLK DW[29] VGND VGND VPWR VPWR
+ REGF\[3\].RFW.BIT\[29\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_12_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_12_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[9\].RFW.BIT\[23\].FF REGF\[9\].RFW.CG\[2\]/GCLK DW[23] VGND VGND VPWR VPWR
+ REGF\[9\].RFW.BIT\[23\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_12_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[15\].RFW.BIT\[13\].FF REGF\[15\].RFW.CG\[1\]/GCLK DW[13] VGND VGND VPWR VPWR
+ REGF\[15\].RFW.BIT\[13\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[18\].RFW.BIT\[11\].OBUF1 REGF\[18\].RFW.BIT\[11\].FF/Q REGF\[18\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[11] sky130_fd_sc_hd__ebufn_2
XREGF\[31\].RFW.BIT\[16\].FF REGF\[31\].RFW.CG\[2\]/GCLK DW[16] VGND VGND VPWR VPWR
+ REGF\[31\].RFW.BIT\[16\].FF/Q sky130_fd_sc_hd__dfxtp_1
XDEC1.D2.AND6 DEC1.D2.AND7/A DEC1.D2.AND7/B DEC1.D2.AND7/C DEC1.D2.AND7/D VGND VGND
+ VPWR VPWR DEC1.D2.AND6/X sky130_fd_sc_hd__and4b_2
XREGF\[14\].RFW.INV2\[3\] DEC1.D1.AND6/X VGND VGND VPWR VPWR REGF\[14\].RFW.INV2\[3\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_37_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_37_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_24_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_37_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_17_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[19\].RFW.BIT\[27\].OBUF2 REGF\[19\].RFW.BIT\[27\].FF/Q REGF\[19\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[27] sky130_fd_sc_hd__ebufn_2
Xfill_53_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_53_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[28\].RFW.BIT\[7\].OBUF2 REGF\[28\].RFW.BIT\[7\].FF/Q REGF\[28\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[7] sky130_fd_sc_hd__ebufn_2
XREGF\[11\].RFW.BIT\[29\].OBUF1 REGF\[11\].RFW.BIT\[29\].FF/Q REGF\[11\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[29] sky130_fd_sc_hd__ebufn_2
XREGF\[20\].RFW.BIT\[29\].FF REGF\[20\].RFW.CG\[3\]/GCLK DW[29] VGND VGND VPWR VPWR
+ REGF\[20\].RFW.BIT\[29\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[23\].RFW.BIT\[1\].OBUF1 REGF\[23\].RFW.BIT\[1\].FF/Q REGF\[23\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[1] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.BIT\[16\].OBUF2 REGF\[24\].RFW.BIT\[16\].FF/Q REGF\[24\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[16] sky130_fd_sc_hd__ebufn_2
Xfill_9_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_9_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_9_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_9_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC2.D.AND0 RW[3] RW[4] DEC2.TIE/HI VGND VGND VPWR VPWR DEC2.D.AND0/Y sky130_fd_sc_hd__nor3b_4
Xfill_9_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[26\].RFW.BIT\[23\].FF REGF\[26\].RFW.CG\[2\]/GCLK DW[23] VGND VGND VPWR VPWR
+ REGF\[26\].RFW.BIT\[23\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[2\].RFW.BIT\[21\].OBUF1 REGF\[2\].RFW.BIT\[21\].FF/Q REGF\[2\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[21] sky130_fd_sc_hd__ebufn_2
Xfill_50_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[14\].RFW.BIT\[14\].OBUF1 REGF\[14\].RFW.BIT\[14\].FF/Q REGF\[14\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[14] sky130_fd_sc_hd__ebufn_2
Xfill_43_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[7\].RFW.INV1\[0\] DEC0.D0.AND7/X VGND VGND VPWR VPWR REGF\[7\].RFW.INV1\[0\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_36_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[21\].RFW.BIT\[5\].OBUF2 REGF\[21\].RFW.BIT\[5\].FF/Q REGF\[21\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[5] sky130_fd_sc_hd__ebufn_2
Xtap_10_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_58_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[19\].OBUF2 REGF\[20\].RFW.BIT\[19\].FF/Q REGF\[20\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[19] sky130_fd_sc_hd__ebufn_2
Xfill_58_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_58_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_58_17 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.BIT\[22\].OBUF2 REGF\[6\].RFW.BIT\[22\].FF/Q REGF\[6\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[22] sky130_fd_sc_hd__ebufn_2
Xtap_1_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[25\].RFW.BIT\[1\].OBUF1 REGF\[25\].RFW.BIT\[1\].FF/Q REGF\[25\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[1] sky130_fd_sc_hd__ebufn_2
XREGF\[18\].RFW.BIT\[15\].OBUF2 REGF\[18\].RFW.BIT\[15\].FF/Q REGF\[18\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[15] sky130_fd_sc_hd__ebufn_2
XREGF\[10\].RFW.BIT\[17\].OBUF1 REGF\[10\].RFW.BIT\[17\].FF/Q REGF\[10\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[17] sky130_fd_sc_hd__ebufn_2
XREGF\[11\].RFW.BIT\[30\].OBUF1 REGF\[11\].RFW.BIT\[30\].FF/Q REGF\[11\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[30] sky130_fd_sc_hd__ebufn_2
Xfill_23_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_23_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_23_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_23_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XREGF\[23\].RFW.BIT\[5\].OBUF2 REGF\[23\].RFW.BIT\[5\].FF/Q REGF\[23\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[5] sky130_fd_sc_hd__ebufn_2
Xfill_22_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_15_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[2\].RFW.BIT\[25\].OBUF2 REGF\[2\].RFW.BIT\[25\].FF/Q REGF\[2\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[25] sky130_fd_sc_hd__ebufn_2
XREGF\[25\].RFW.CGAND DEC2.D3.AND1/X WE VGND VGND VPWR VPWR REGF\[25\].RFW.CGAND/X
+ sky130_fd_sc_hd__and2_1
XREGF\[14\].RFW.BIT\[18\].OBUF2 REGF\[14\].RFW.BIT\[18\].FF/Q REGF\[14\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[18] sky130_fd_sc_hd__ebufn_2
XREGF\[15\].RFW.BIT\[31\].OBUF2 REGF\[15\].RFW.BIT\[31\].FF/Q REGF\[15\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[31] sky130_fd_sc_hd__ebufn_2
XREGF\[16\].RFW.BIT\[19\].FF REGF\[16\].RFW.CG\[2\]/GCLK DW[19] VGND VGND VPWR VPWR
+ REGF\[16\].RFW.BIT\[19\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[6\].RFW.BIT\[31\].FF REGF\[6\].RFW.CG\[3\]/GCLK DW[31] VGND VGND VPWR VPWR
+ REGF\[6\].RFW.BIT\[31\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[12\].RFW.BIT\[21\].FF REGF\[12\].RFW.CG\[2\]/GCLK DW[21] VGND VGND VPWR VPWR
+ REGF\[12\].RFW.BIT\[21\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[20\].RFW.BIT\[20\].OBUF2 REGF\[20\].RFW.BIT\[20\].FF/Q REGF\[20\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[20] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[1\].OBUF1 REGF\[27\].RFW.BIT\[1\].FF/Q REGF\[27\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[1] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[10\].OBUF2 REGF\[5\].RFW.BIT\[10\].FF/Q REGF\[5\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[10] sky130_fd_sc_hd__ebufn_2
XREGF\[1\].RFW.INV2\[1\] DEC1.D0.AND1/X VGND VGND VPWR VPWR REGF\[1\].RFW.INV2\[1\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_44_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_60_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xtap_56_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[25\].RFW.BIT\[5\].OBUF2 REGF\[25\].RFW.BIT\[5\].FF/Q REGF\[25\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[5] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[29\].FF REGF\[27\].RFW.CG\[3\]/GCLK DW[29] VGND VGND VPWR VPWR
+ REGF\[27\].RFW.BIT\[29\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_49_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[23\].RFW.BIT\[31\].FF REGF\[23\].RFW.CG\[3\]/GCLK DW[31] VGND VGND VPWR VPWR
+ REGF\[23\].RFW.BIT\[31\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_18_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_18_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_34_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[1\].RFW.BIT\[13\].OBUF2 REGF\[1\].RFW.BIT\[13\].FF/Q REGF\[1\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[13] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.BIT\[1\].OBUF1 REGF\[29\].RFW.BIT\[1\].FF/Q REGF\[29\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[1] sky130_fd_sc_hd__ebufn_2
Xfill_50_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XDEC2.D0.ABUF\[1\] RW[1] VGND VGND VPWR VPWR DEC2.D0.AND7/B sky130_fd_sc_hd__clkbuf_2
XREGF\[7\].RFW.BIT\[14\].FF REGF\[7\].RFW.CG\[1\]/GCLK DW[14] VGND VGND VPWR VPWR
+ REGF\[7\].RFW.BIT\[14\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_6_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_6_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_59_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_6_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[30\].RFW.CG\[2\] CLK REGF\[30\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[30\].RFW.CG\[2\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_20_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[29\].RFW.BIT\[16\].OBUF1 REGF\[29\].RFW.BIT\[16\].FF/Q REGF\[29\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[16] sky130_fd_sc_hd__ebufn_2
Xfill_13_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XREGF\[27\].RFW.BIT\[5\].OBUF2 REGF\[27\].RFW.BIT\[5\].FF/Q REGF\[27\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[5] sky130_fd_sc_hd__ebufn_2
XREGF\[10\].RFW.BIT\[22\].OBUF2 REGF\[10\].RFW.BIT\[22\].FF/Q REGF\[10\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[22] sky130_fd_sc_hd__ebufn_2
Xtap_28_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[24\].RFW.BIT\[14\].FF REGF\[24\].RFW.CG\[1\]/GCLK DW[14] VGND VGND VPWR VPWR
+ REGF\[24\].RFW.BIT\[14\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_39_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_16_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_55_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_55_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[20\].RFW.BIT\[3\].OBUF2 REGF\[20\].RFW.BIT\[3\].FF/Q REGF\[20\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[3] sky130_fd_sc_hd__ebufn_2
Xtap_32_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_61_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[25\].RFW.BIT\[19\].OBUF1 REGF\[25\].RFW.BIT\[19\].FF/Q REGF\[25\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[19] sky130_fd_sc_hd__ebufn_2
Xtap_54_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[13\].RFW.BIT\[27\].FF REGF\[13\].RFW.CG\[3\]/GCLK DW[27] VGND VGND VPWR VPWR
+ REGF\[13\].RFW.BIT\[27\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[16\].RFW.INV2\[0\] DEC1.D2.AND0/Y VGND VGND VPWR VPWR REGF\[16\].RFW.INV2\[0\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_20_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_47_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_20_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_20_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.BIT\[21\].OBUF1 REGF\[31\].RFW.BIT\[21\].FF/Q REGF\[31\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[21] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.BIT\[21\].FF REGF\[19\].RFW.CG\[2\]/GCLK DW[21] VGND VGND VPWR VPWR
+ REGF\[19\].RFW.BIT\[21\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_29_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_29_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_29_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_29_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[29\].RFW.BIT\[5\].OBUF2 REGF\[29\].RFW.BIT\[5\].FF/Q REGF\[29\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[5] sky130_fd_sc_hd__ebufn_2
Xfill_45_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_45_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_45_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[31\].RFW.BIT\[8\].OBUF1 REGF\[31\].RFW.BIT\[8\].FF/Q REGF\[31\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[8] sky130_fd_sc_hd__ebufn_2
Xfill_61_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_61_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[7\].RFW.CG\[2\] CLK REGF\[7\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[7\].RFW.CG\[2\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[22\].RFW.BIT\[3\].OBUF2 REGF\[22\].RFW.BIT\[3\].FF/Q REGF\[22\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[3] sky130_fd_sc_hd__ebufn_2
XREGF\[7\].RFW.BIT\[25\].OBUF1 REGF\[7\].RFW.BIT\[25\].FF/Q REGF\[7\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[25] sky130_fd_sc_hd__ebufn_2
Xfill_9_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[19\].RFW.BIT\[18\].OBUF1 REGF\[19\].RFW.BIT\[18\].FF/Q REGF\[19\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[18] sky130_fd_sc_hd__ebufn_2
XREGF\[12\].RFW.INV1\[1\] DEC0.D1.AND4/X VGND VGND VPWR VPWR REGF\[12\].RFW.INV1\[1\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[25\].RFW.BIT\[20\].OBUF1 REGF\[25\].RFW.BIT\[20\].FF/Q REGF\[25\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[20] sky130_fd_sc_hd__ebufn_2
XREGF\[28\].RFW.INV1\[2\] DEC0.D3.AND4/X VGND VGND VPWR VPWR REGF\[28\].RFW.INV1\[2\]/Y
+ sky130_fd_sc_hd__inv_4
Xtap_40_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[4\].RFW.BIT\[22\].FF REGF\[4\].RFW.CG\[2\]/GCLK DW[22] VGND VGND VPWR VPWR
+ REGF\[4\].RFW.BIT\[22\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[10\].RFW.BIT\[12\].FF REGF\[10\].RFW.CG\[1\]/GCLK DW[12] VGND VGND VPWR VPWR
+ REGF\[10\].RFW.BIT\[12\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_19_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.BIT\[25\].OBUF2 REGF\[31\].RFW.BIT\[25\].FF/Q REGF\[31\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[25] sky130_fd_sc_hd__ebufn_2
Xfill_15_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_15_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_15_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC0.D1.ENBUF DEC0.D.AND1/X VGND VGND VPWR VPWR DEC0.D1.AND7/D sky130_fd_sc_hd__clkbuf_2
Xfill_15_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_15_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_31_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[24\].RFW.BIT\[3\].OBUF2 REGF\[24\].RFW.BIT\[3\].FF/Q REGF\[24\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[3] sky130_fd_sc_hd__ebufn_2
XREGF\[3\].RFW.BIT\[28\].OBUF1 REGF\[3\].RFW.BIT\[28\].FF/Q REGF\[3\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[28] sky130_fd_sc_hd__ebufn_2
Xfill_31_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_31_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_31_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XREGF\[29\].RFW.BIT\[21\].OBUF2 REGF\[29\].RFW.BIT\[21\].FF/Q REGF\[29\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[21] sky130_fd_sc_hd__ebufn_2
XREGF\[19\].RFW.BIT\[5\].FF REGF\[19\].RFW.CG\[0\]/GCLK DW[5] VGND VGND VPWR VPWR
+ REGF\[19\].RFW.BIT\[5\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[21\].RFW.BIT\[23\].OBUF1 REGF\[21\].RFW.BIT\[23\].FF/Q REGF\[21\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[23] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.BIT\[22\].FF REGF\[21\].RFW.CG\[2\]/GCLK DW[22] VGND VGND VPWR VPWR
+ REGF\[21\].RFW.BIT\[22\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_54_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_47_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[6\].RFW.BIT\[13\].OBUF1 REGF\[6\].RFW.BIT\[13\].FF/Q REGF\[6\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[13] sky130_fd_sc_hd__ebufn_2
Xfill_3_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_3_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_3_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XDEC1.D1.ABUF\[2\] RB[2] VGND VGND VPWR VPWR DEC1.D1.AND7/C sky130_fd_sc_hd__clkbuf_2
Xfill_3_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_2_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.BIT\[7\].FF REGF\[18\].RFW.CG\[0\]/GCLK DW[7] VGND VGND VPWR VPWR
+ REGF\[18\].RFW.BIT\[7\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[7\].RFW.BIT\[29\].OBUF2 REGF\[7\].RFW.BIT\[29\].FF/Q REGF\[7\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[29] sky130_fd_sc_hd__ebufn_2
XREGF\[25\].RFW.BIT\[24\].OBUF2 REGF\[25\].RFW.BIT\[24\].FF/Q REGF\[25\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[24] sky130_fd_sc_hd__ebufn_2
XREGF\[17\].RFW.BIT\[9\].FF REGF\[17\].RFW.CG\[1\]/GCLK DW[9] VGND VGND VPWR VPWR
+ REGF\[17\].RFW.BIT\[9\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[30\].RFW.BIT\[13\].OBUF2 REGF\[30\].RFW.BIT\[13\].FF/Q REGF\[30\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[13] sky130_fd_sc_hd__ebufn_2
XREGF\[26\].RFW.BIT\[3\].OBUF2 REGF\[26\].RFW.BIT\[3\].FF/Q REGF\[26\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[3] sky130_fd_sc_hd__ebufn_2
Xfill_52_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[2\].RFW.BIT\[16\].OBUF1 REGF\[2\].RFW.BIT\[16\].FF/Q REGF\[2\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[16] sky130_fd_sc_hd__ebufn_2
XREGF\[15\].RFW.BIT\[22\].OBUF1 REGF\[15\].RFW.BIT\[22\].FF/Q REGF\[15\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[22] sky130_fd_sc_hd__ebufn_2
XREGF\[22\].RFW.INV2\[3\] DEC1.D2.AND6/X VGND VGND VPWR VPWR REGF\[22\].RFW.INV2\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[20\].RFW.BIT\[11\].OBUF1 REGF\[20\].RFW.BIT\[11\].FF/Q REGF\[20\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[11] sky130_fd_sc_hd__ebufn_2
Xtap_31_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_38_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgenblk1.RFW0.INV2\[1\] DEC1.D0.AND0/Y VGND VGND VPWR VPWR genblk1.RFW0.INV2\[1\]/Y
+ sky130_fd_sc_hd__inv_4
Xtap_24_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_26_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_26_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[21\].RFW.BIT\[27\].OBUF2 REGF\[21\].RFW.BIT\[27\].FF/Q REGF\[21\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[27] sky130_fd_sc_hd__ebufn_2
Xfill_42_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_42_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[7\].RFW.BIT\[30\].OBUF2 REGF\[7\].RFW.BIT\[30\].FF/Q REGF\[7\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[30] sky130_fd_sc_hd__ebufn_2
XREGF\[6\].RFW.BIT\[17\].OBUF2 REGF\[6\].RFW.BIT\[17\].FF/Q REGF\[6\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[17] sky130_fd_sc_hd__ebufn_2
XREGF\[5\].RFW.BIT\[28\].FF REGF\[5\].RFW.CG\[3\]/GCLK DW[28] VGND VGND VPWR VPWR
+ REGF\[5\].RFW.BIT\[28\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[19\].RFW.BIT\[23\].OBUF2 REGF\[19\].RFW.BIT\[23\].FF/Q REGF\[19\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[23] sky130_fd_sc_hd__ebufn_2
XREGF\[11\].RFW.BIT\[18\].FF REGF\[11\].RFW.CG\[2\]/GCLK DW[18] VGND VGND VPWR VPWR
+ REGF\[11\].RFW.BIT\[18\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[28\].RFW.BIT\[3\].OBUF2 REGF\[28\].RFW.BIT\[3\].FF/Q REGF\[28\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[3] sky130_fd_sc_hd__ebufn_2
Xfill_52_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[1\].RFW.BIT\[30\].FF REGF\[1\].RFW.CG\[3\]/GCLK DW[30] VGND VGND VPWR VPWR
+ REGF\[1\].RFW.BIT\[30\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[24\].RFW.BIT\[12\].OBUF2 REGF\[24\].RFW.BIT\[12\].FF/Q REGF\[24\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[12] sky130_fd_sc_hd__ebufn_2
XREGF\[11\].RFW.BIT\[25\].OBUF1 REGF\[11\].RFW.BIT\[25\].FF/Q REGF\[11\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[25] sky130_fd_sc_hd__ebufn_2
Xfill_45_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[17\].RFW.BIT\[12\].FF REGF\[17\].RFW.CG\[1\]/GCLK DW[12] VGND VGND VPWR VPWR
+ REGF\[17\].RFW.BIT\[12\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_38_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_0_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[30\].RFW.BIT\[6\].OBUF1 REGF\[30\].RFW.BIT\[6\].FF/Q REGF\[30\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[6] sky130_fd_sc_hd__ebufn_2
XDEC2.D1.AND5 DEC2.D1.AND7/B DEC2.D1.AND7/A DEC2.D1.AND7/C DEC2.D1.AND7/D VGND VGND
+ VPWR VPWR DEC2.D1.AND5/X sky130_fd_sc_hd__and4b_2
XREGF\[14\].RFW.BIT\[10\].OBUF1 REGF\[14\].RFW.BIT\[10\].FF/Q REGF\[14\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[10] sky130_fd_sc_hd__ebufn_2
XREGF\[21\].RFW.BIT\[1\].OBUF2 REGF\[21\].RFW.BIT\[1\].FF/Q REGF\[21\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[1] sky130_fd_sc_hd__ebufn_2
XREGF\[22\].RFW.BIT\[28\].FF REGF\[22\].RFW.CG\[3\]/GCLK DW[28] VGND VGND VPWR VPWR
+ REGF\[22\].RFW.BIT\[28\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_10_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_47_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[28\].RFW.BIT\[22\].FF REGF\[28\].RFW.CG\[2\]/GCLK DW[22] VGND VGND VPWR VPWR
+ REGF\[28\].RFW.BIT\[22\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[15\].RFW.BIT\[26\].OBUF2 REGF\[15\].RFW.BIT\[26\].FF/Q REGF\[15\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[26] sky130_fd_sc_hd__ebufn_2
Xtap_24_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[15\].OBUF2 REGF\[20\].RFW.BIT\[15\].FF/Q REGF\[20\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[15] sky130_fd_sc_hd__ebufn_2
Xtap_40_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_12_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_12_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_12_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.BIT\[11\].OBUF2 REGF\[18\].RFW.BIT\[11\].FF/Q REGF\[18\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[11] sky130_fd_sc_hd__ebufn_2
XREGF\[10\].RFW.BIT\[13\].OBUF1 REGF\[10\].RFW.BIT\[13\].FF/Q REGF\[10\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[13] sky130_fd_sc_hd__ebufn_2
XREGF\[2\].RFW.BIT\[13\].FF REGF\[2\].RFW.CG\[1\]/GCLK DW[13] VGND VGND VPWR VPWR
+ REGF\[2\].RFW.BIT\[13\].FF/Q sky130_fd_sc_hd__dfxtp_1
XDEC1.D2.AND7 DEC1.D2.AND7/A DEC1.D2.AND7/B DEC1.D2.AND7/C DEC1.D2.AND7/D VGND VGND
+ VPWR VPWR DEC1.D2.AND7/X sky130_fd_sc_hd__and4_2
Xfill_37_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_37_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_37_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_37_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_17_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_0_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_53_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_53_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_53_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[11\].RFW.BIT\[29\].OBUF2 REGF\[11\].RFW.BIT\[29\].FF/Q REGF\[11\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[29] sky130_fd_sc_hd__ebufn_2
XREGF\[23\].RFW.BIT\[1\].OBUF2 REGF\[23\].RFW.BIT\[1\].FF/Q REGF\[23\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[1] sky130_fd_sc_hd__ebufn_2
XREGF\[24\].RFW.CGAND DEC2.D3.AND0/Y WE VGND VGND VPWR VPWR REGF\[24\].RFW.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_9_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_9_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_9_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC2.D.AND1 RW[4] RW[3] DEC2.TIE/HI VGND VGND VPWR VPWR DEC2.D.AND1/X sky130_fd_sc_hd__and3b_4
Xfill_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_9_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[2\].RFW.BIT\[21\].OBUF2 REGF\[2\].RFW.BIT\[21\].FF/Q REGF\[2\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[21] sky130_fd_sc_hd__ebufn_2
Xfill_50_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_43_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[14\].RFW.BIT\[14\].OBUF2 REGF\[14\].RFW.BIT\[14\].FF/Q REGF\[14\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[14] sky130_fd_sc_hd__ebufn_2
Xfill_36_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_29_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_58_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_58_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[18\].RFW.BIT\[18\].FF REGF\[18\].RFW.CG\[2\]/GCLK DW[18] VGND VGND VPWR VPWR
+ REGF\[18\].RFW.BIT\[18\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[8\].RFW.BIT\[30\].FF REGF\[8\].RFW.CG\[3\]/GCLK DW[30] VGND VGND VPWR VPWR
+ REGF\[8\].RFW.BIT\[30\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[14\].RFW.BIT\[20\].FF REGF\[14\].RFW.CG\[2\]/GCLK DW[20] VGND VGND VPWR VPWR
+ REGF\[14\].RFW.BIT\[20\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_1_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[25\].RFW.BIT\[1\].OBUF2 REGF\[25\].RFW.BIT\[1\].FF/Q REGF\[25\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[1] sky130_fd_sc_hd__ebufn_2
XREGF\[30\].RFW.BIT\[23\].FF REGF\[30\].RFW.CG\[2\]/GCLK DW[23] VGND VGND VPWR VPWR
+ REGF\[30\].RFW.BIT\[23\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[11\].RFW.BIT\[30\].OBUF2 REGF\[11\].RFW.BIT\[30\].FF/Q REGF\[11\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[30] sky130_fd_sc_hd__ebufn_2
XREGF\[10\].RFW.BIT\[17\].OBUF2 REGF\[10\].RFW.BIT\[17\].FF/Q REGF\[10\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[17] sky130_fd_sc_hd__ebufn_2
Xfill_23_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_23_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_23_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_23_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_23_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[29\].RFW.BIT\[28\].FF REGF\[29\].RFW.CG\[3\]/GCLK DW[28] VGND VGND VPWR VPWR
+ REGF\[29\].RFW.BIT\[28\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_48_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[26\].RFW.BIT\[27\].OBUF1 REGF\[26\].RFW.BIT\[27\].FF/Q REGF\[26\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[27] sky130_fd_sc_hd__ebufn_2
XREGF\[25\].RFW.BIT\[30\].FF REGF\[25\].RFW.CG\[3\]/GCLK DW[30] VGND VGND VPWR VPWR
+ REGF\[25\].RFW.BIT\[30\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_22_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_15_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.BIT\[16\].OBUF1 REGF\[31\].RFW.BIT\[16\].FF/Q REGF\[31\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[16] sky130_fd_sc_hd__ebufn_2
XREGF\[4\].RFW.INV2\[2\] DEC1.D0.AND4/X VGND VGND VPWR VPWR REGF\[4\].RFW.INV2\[2\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[29\].RFW.BIT\[12\].OBUF1 REGF\[29\].RFW.BIT\[12\].FF/Q REGF\[29\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[12] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[1\].OBUF2 REGF\[27\].RFW.BIT\[1\].FF/Q REGF\[27\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[1] sky130_fd_sc_hd__ebufn_2
XREGF\[3\].RFW.BIT\[19\].FF REGF\[3\].RFW.CG\[2\]/GCLK DW[19] VGND VGND VPWR VPWR
+ REGF\[3\].RFW.BIT\[19\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[15\].RFW.BIT\[0\].FF REGF\[15\].RFW.CG\[0\]/GCLK DW[0] VGND VGND VPWR VPWR
+ REGF\[15\].RFW.BIT\[0\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[9\].RFW.BIT\[13\].FF REGF\[9\].RFW.CG\[1\]/GCLK DW[13] VGND VGND VPWR VPWR
+ REGF\[9\].RFW.BIT\[13\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[24\].RFW.INV2\[0\] DEC1.D3.AND0/Y VGND VGND VPWR VPWR REGF\[24\].RFW.INV2\[0\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_60_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_56_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[14\].RFW.BIT\[2\].FF REGF\[14\].RFW.CG\[0\]/GCLK DW[2] VGND VGND VPWR VPWR
+ REGF\[14\].RFW.BIT\[2\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_46_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_18_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[20\].RFW.BIT\[19\].FF REGF\[20\].RFW.CG\[2\]/GCLK DW[19] VGND VGND VPWR VPWR
+ REGF\[20\].RFW.BIT\[19\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[25\].RFW.BIT\[15\].OBUF1 REGF\[25\].RFW.BIT\[15\].FF/Q REGF\[25\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[15] sky130_fd_sc_hd__ebufn_2
Xfill_18_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_18_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[26\].RFW.BIT\[13\].FF REGF\[26\].RFW.CG\[1\]/GCLK DW[13] VGND VGND VPWR VPWR
+ REGF\[26\].RFW.BIT\[13\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_34_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_34_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[13\].RFW.BIT\[4\].FF REGF\[13\].RFW.CG\[0\]/GCLK DW[4] VGND VGND VPWR VPWR
+ REGF\[13\].RFW.BIT\[4\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[29\].RFW.BIT\[1\].OBUF2 REGF\[29\].RFW.BIT\[1\].FF/Q REGF\[29\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[1] sky130_fd_sc_hd__ebufn_2
XREGF\[3\].RFW.CG\[1\] CLK REGF\[3\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[3\].RFW.CG\[1\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
Xfill_50_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfill_50_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_6_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_6_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.BIT\[4\].OBUF1 REGF\[31\].RFW.BIT\[4\].FF/Q REGF\[31\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[4] sky130_fd_sc_hd__ebufn_2
Xfill_59_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_59_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_6_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[28\].RFW.BIT\[0\].FF REGF\[28\].RFW.CG\[0\]/GCLK DW[0] VGND VGND VPWR VPWR
+ REGF\[28\].RFW.BIT\[0\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[15\].RFW.BIT\[26\].FF REGF\[15\].RFW.CG\[3\]/GCLK DW[26] VGND VGND VPWR VPWR
+ REGF\[15\].RFW.BIT\[26\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[12\].RFW.BIT\[6\].FF REGF\[12\].RFW.CG\[0\]/GCLK DW[6] VGND VGND VPWR VPWR
+ REGF\[12\].RFW.BIT\[6\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[31\].RFW.BIT\[29\].FF REGF\[31\].RFW.CG\[3\]/GCLK DW[29] VGND VGND VPWR VPWR
+ REGF\[31\].RFW.BIT\[29\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_20_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[20\].RFW.INV1\[1\] DEC0.D2.AND4/X VGND VGND VPWR VPWR REGF\[20\].RFW.INV1\[1\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[16\].RFW.BIT\[29\].OBUF1 REGF\[16\].RFW.BIT\[29\].FF/Q REGF\[16\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[29] sky130_fd_sc_hd__ebufn_2
XREGF\[29\].RFW.CG\[0\] CLK REGF\[29\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[29\].RFW.CG\[0\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[29\].RFW.BIT\[16\].OBUF2 REGF\[29\].RFW.BIT\[16\].FF/Q REGF\[29\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[16] sky130_fd_sc_hd__ebufn_2
Xfill_13_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[21\].RFW.BIT\[18\].OBUF1 REGF\[21\].RFW.BIT\[18\].FF/Q REGF\[21\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[18] sky130_fd_sc_hd__ebufn_2
XREGF\[22\].RFW.BIT\[31\].OBUF1 REGF\[22\].RFW.BIT\[31\].FF/Q REGF\[22\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[31] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[2\].FF REGF\[27\].RFW.CG\[0\]/GCLK DW[2] VGND VGND VPWR VPWR
+ REGF\[27\].RFW.BIT\[2\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[7\].RFW.BIT\[21\].OBUF1 REGF\[7\].RFW.BIT\[21\].FF/Q REGF\[7\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[21] sky130_fd_sc_hd__ebufn_2
XREGF\[11\].RFW.BIT\[8\].FF REGF\[11\].RFW.CG\[1\]/GCLK DW[8] VGND VGND VPWR VPWR
+ REGF\[11\].RFW.BIT\[8\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[19\].RFW.BIT\[14\].OBUF1 REGF\[19\].RFW.BIT\[14\].FF/Q REGF\[19\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[14] sky130_fd_sc_hd__ebufn_2
Xtap_28_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[19\].RFW.INV2\[1\] DEC1.D2.AND3/X VGND VGND VPWR VPWR REGF\[19\].RFW.INV2\[1\]/Y
+ sky130_fd_sc_hd__inv_4
Xfill_55_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_32_12 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[26\].RFW.BIT\[4\].FF REGF\[26\].RFW.CG\[0\]/GCLK DW[4] VGND VGND VPWR VPWR
+ REGF\[26\].RFW.BIT\[4\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xtap_61_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_54_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[18\].RFW.CG\[3\] CLK REGF\[18\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[18\].RFW.CG\[3\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[25\].RFW.BIT\[19\].OBUF2 REGF\[25\].RFW.BIT\[19\].FF/Q REGF\[25\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[19] sky130_fd_sc_hd__ebufn_2
Xfill_20_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_20_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_20_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_47_1 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[31\].RFW.BIT\[21\].OBUF2 REGF\[31\].RFW.BIT\[21\].FF/Q REGF\[31\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[21] sky130_fd_sc_hd__ebufn_2
Xfill_29_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_29_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_29_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_29_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XREGF\[25\].RFW.BIT\[6\].FF REGF\[25\].RFW.CG\[0\]/GCLK DW[6] VGND VGND VPWR VPWR
+ REGF\[25\].RFW.BIT\[6\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[3\].RFW.BIT\[24\].OBUF1 REGF\[3\].RFW.BIT\[24\].FF/Q REGF\[3\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[24] sky130_fd_sc_hd__ebufn_2
XREGF\[15\].RFW.BIT\[17\].OBUF1 REGF\[15\].RFW.BIT\[17\].FF/Q REGF\[15\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[17] sky130_fd_sc_hd__ebufn_2
XREGF\[6\].RFW.BIT\[21\].FF REGF\[6\].RFW.CG\[2\]/GCLK DW[21] VGND VGND VPWR VPWR
+ REGF\[6\].RFW.BIT\[21\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[16\].RFW.BIT\[30\].OBUF1 REGF\[16\].RFW.BIT\[30\].FF/Q REGF\[16\].RFW.INV1\[3\]/Y
+ VGND VGND VPWR VPWR DA[30] sky130_fd_sc_hd__ebufn_2
Xfill_45_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_45_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[12\].RFW.BIT\[11\].FF REGF\[12\].RFW.CG\[1\]/GCLK DW[11] VGND VGND VPWR VPWR
+ REGF\[12\].RFW.BIT\[11\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_45_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_45_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[31\].RFW.BIT\[8\].OBUF2 REGF\[31\].RFW.BIT\[8\].FF/Q REGF\[31\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[8] sky130_fd_sc_hd__ebufn_2
Xfill_61_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_61_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_61_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[24\].RFW.BIT\[8\].FF REGF\[24\].RFW.CG\[1\]/GCLK DW[8] VGND VGND VPWR VPWR
+ REGF\[24\].RFW.BIT\[8\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[17\].RFW.CG\[0\] CLK REGF\[17\].RFW.CGAND/X VGND VGND VPWR VPWR REGF\[17\].RFW.CG\[0\]/GCLK
+ sky130_fd_sc_hd__dlclkp_1
XREGF\[15\].RFW.INV1\[2\] DEC0.D1.AND7/X VGND VGND VPWR VPWR REGF\[15\].RFW.INV1\[2\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[7\].RFW.BIT\[25\].OBUF2 REGF\[7\].RFW.BIT\[25\].FF/Q REGF\[7\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[25] sky130_fd_sc_hd__ebufn_2
XREGF\[27\].RFW.BIT\[19\].FF REGF\[27\].RFW.CG\[2\]/GCLK DW[19] VGND VGND VPWR VPWR
+ REGF\[27\].RFW.BIT\[19\].FF/Q sky130_fd_sc_hd__dfxtp_1
Xfill_11_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_9_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[23\].RFW.BIT\[21\].FF REGF\[23\].RFW.CG\[2\]/GCLK DW[21] VGND VGND VPWR VPWR
+ REGF\[23\].RFW.BIT\[21\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[19\].RFW.BIT\[18\].OBUF2 REGF\[19\].RFW.BIT\[18\].FF/Q REGF\[19\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[18] sky130_fd_sc_hd__ebufn_2
XREGF\[30\].RFW.INV2\[3\] DEC1.D3.AND6/X VGND VGND VPWR VPWR REGF\[30\].RFW.INV2\[3\]/Y
+ sky130_fd_sc_hd__inv_4
XREGF\[25\].RFW.BIT\[20\].OBUF2 REGF\[25\].RFW.BIT\[20\].FF/Q REGF\[25\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[20] sky130_fd_sc_hd__ebufn_2
Xtap_40_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_26_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[9\].RFW.BIT\[5\].FF REGF\[9\].RFW.CG\[0\]/GCLK DW[5] VGND VGND VPWR VPWR REGF\[9\].RFW.BIT\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xtap_19_5 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[2\].RFW.BIT\[12\].OBUF1 REGF\[2\].RFW.BIT\[12\].FF/Q REGF\[2\].RFW.INV1\[1\]/Y
+ VGND VGND VPWR VPWR DA[12] sky130_fd_sc_hd__ebufn_2
Xfill_15_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_15_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_15_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_15_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_15_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_31_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XREGF\[3\].RFW.BIT\[28\].OBUF2 REGF\[3\].RFW.BIT\[28\].FF/Q REGF\[3\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[28] sky130_fd_sc_hd__ebufn_2
XREGF\[8\].RFW.BIT\[7\].FF REGF\[8\].RFW.CG\[0\]/GCLK DW[7] VGND VGND VPWR VPWR REGF\[8\].RFW.BIT\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xfill_31_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_31_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_31_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_31_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[21\].RFW.BIT\[23\].OBUF2 REGF\[21\].RFW.BIT\[23\].FF/Q REGF\[21\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[23] sky130_fd_sc_hd__ebufn_2
Xfill_47_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_56_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XREGF\[6\].RFW.BIT\[13\].OBUF2 REGF\[6\].RFW.BIT\[13\].FF/Q REGF\[6\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[13] sky130_fd_sc_hd__ebufn_2
Xfill_3_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfill_3_13 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_3_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[7\].RFW.BIT\[9\].FF REGF\[7\].RFW.CG\[1\]/GCLK DW[9] VGND VGND VPWR VPWR REGF\[7\].RFW.BIT\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
Xfill_2_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[11\].RFW.BIT\[21\].OBUF1 REGF\[11\].RFW.BIT\[21\].FF/Q REGF\[11\].RFW.INV1\[2\]/Y
+ VGND VGND VPWR VPWR DA[21] sky130_fd_sc_hd__ebufn_2
XREGF\[30\].RFW.BIT\[2\].OBUF1 REGF\[30\].RFW.BIT\[2\].FF/Q REGF\[30\].RFW.INV1\[0\]/Y
+ VGND VGND VPWR VPWR DA[2] sky130_fd_sc_hd__ebufn_2
Xfill_59_0 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[7\].RFW.BIT\[27\].FF REGF\[7\].RFW.CG\[3\]/GCLK DW[27] VGND VGND VPWR VPWR
+ REGF\[7\].RFW.BIT\[27\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[13\].RFW.BIT\[17\].FF REGF\[13\].RFW.CG\[2\]/GCLK DW[17] VGND VGND VPWR VPWR
+ REGF\[13\].RFW.BIT\[17\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[19\].RFW.BIT\[11\].FF REGF\[19\].RFW.CG\[1\]/GCLK DW[11] VGND VGND VPWR VPWR
+ REGF\[19\].RFW.BIT\[11\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[2\].RFW.BIT\[16\].OBUF2 REGF\[2\].RFW.BIT\[16\].FF/Q REGF\[2\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[16] sky130_fd_sc_hd__ebufn_2
XREGF\[15\].RFW.BIT\[22\].OBUF2 REGF\[15\].RFW.BIT\[22\].FF/Q REGF\[15\].RFW.INV2\[2\]/Y
+ VGND VGND VPWR VPWR DB[22] sky130_fd_sc_hd__ebufn_2
XREGF\[20\].RFW.BIT\[11\].OBUF2 REGF\[20\].RFW.BIT\[11\].FF/Q REGF\[20\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[11] sky130_fd_sc_hd__ebufn_2
Xtap_31_4 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_38_11 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_24_3 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtap_17_2 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[2\].RFW.INV1\[0\] DEC0.D0.AND2/X VGND VGND VPWR VPWR REGF\[2\].RFW.INV1\[0\]/Y
+ sky130_fd_sc_hd__inv_4
Xtap_54_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_26_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_26_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_26_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XREGF\[24\].RFW.BIT\[27\].FF REGF\[24\].RFW.CG\[3\]/GCLK DW[27] VGND VGND VPWR VPWR
+ REGF\[24\].RFW.BIT\[27\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[23\].RFW.CGAND DEC2.D2.AND7/X WE VGND VGND VPWR VPWR REGF\[23\].RFW.CGAND/X
+ sky130_fd_sc_hd__and2_1
Xfill_42_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_42_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfill_52_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XREGF\[11\].RFW.BIT\[25\].OBUF2 REGF\[11\].RFW.BIT\[25\].FF/Q REGF\[11\].RFW.INV2\[3\]/Y
+ VGND VGND VPWR VPWR DB[25] sky130_fd_sc_hd__ebufn_2
Xfill_45_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfill_38_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xfill_0_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XREGF\[30\].RFW.BIT\[6\].OBUF2 REGF\[30\].RFW.BIT\[6\].FF/Q REGF\[30\].RFW.INV2\[0\]/Y
+ VGND VGND VPWR VPWR DB[6] sky130_fd_sc_hd__ebufn_2
XDEC2.D1.AND6 DEC2.D1.AND7/A DEC2.D1.AND7/B DEC2.D1.AND7/C DEC2.D1.AND7/D VGND VGND
+ VPWR VPWR DEC2.D1.AND6/X sky130_fd_sc_hd__and4b_2
XREGF\[4\].RFW.BIT\[12\].FF REGF\[4\].RFW.CG\[1\]/GCLK DW[12] VGND VGND VPWR VPWR
+ REGF\[4\].RFW.BIT\[12\].FF/Q sky130_fd_sc_hd__dfxtp_1
XREGF\[14\].RFW.BIT\[10\].OBUF2 REGF\[14\].RFW.BIT\[10\].FF/Q REGF\[14\].RFW.INV2\[1\]/Y
+ VGND VGND VPWR VPWR DB[10] sky130_fd_sc_hd__ebufn_2
Xtap_10_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XDEC0.D0.ENBUF DEC0.D.AND0/Y VGND VGND VPWR VPWR DEC0.D0.AND7/D sky130_fd_sc_hd__clkbuf_2
.ends

