VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DFFRF_2R1W
  CLASS BLOCK ;
  FOREIGN DFFRF_2R1W ;
  ORIGIN 0.000 0.000 ;
  SIZE 358.800 BY 176.800 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 2.000 ;
    END
  END CLK
  PIN DA[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 2.000 ;
    END
  END DA[0]
  PIN DA[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 2.000 ;
    END
  END DA[10]
  PIN DA[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 2.000 ;
    END
  END DA[11]
  PIN DA[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 2.000 ;
    END
  END DA[12]
  PIN DA[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 2.000 ;
    END
  END DA[13]
  PIN DA[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 2.000 ;
    END
  END DA[14]
  PIN DA[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 2.000 ;
    END
  END DA[15]
  PIN DA[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 2.000 ;
    END
  END DA[16]
  PIN DA[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 2.000 ;
    END
  END DA[17]
  PIN DA[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 2.000 ;
    END
  END DA[18]
  PIN DA[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 2.000 ;
    END
  END DA[19]
  PIN DA[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 2.000 ;
    END
  END DA[1]
  PIN DA[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 2.000 ;
    END
  END DA[20]
  PIN DA[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 2.000 ;
    END
  END DA[21]
  PIN DA[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 2.000 ;
    END
  END DA[22]
  PIN DA[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 0.000 118.590 2.000 ;
    END
  END DA[23]
  PIN DA[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 2.000 ;
    END
  END DA[24]
  PIN DA[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 0.000 128.710 2.000 ;
    END
  END DA[25]
  PIN DA[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 2.000 ;
    END
  END DA[26]
  PIN DA[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 2.000 ;
    END
  END DA[27]
  PIN DA[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 2.000 ;
    END
  END DA[28]
  PIN DA[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.670 0.000 148.950 2.000 ;
    END
  END DA[29]
  PIN DA[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 2.000 ;
    END
  END DA[2]
  PIN DA[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 0.000 154.010 2.000 ;
    END
  END DA[30]
  PIN DA[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 0.000 159.070 2.000 ;
    END
  END DA[31]
  PIN DA[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 2.000 ;
    END
  END DA[3]
  PIN DA[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 2.000 ;
    END
  END DA[4]
  PIN DA[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 0.000 27.510 2.000 ;
    END
  END DA[5]
  PIN DA[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 2.000 ;
    END
  END DA[6]
  PIN DA[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 2.000 ;
    END
  END DA[7]
  PIN DA[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 2.000 ;
    END
  END DA[8]
  PIN DA[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 0.000 47.750 2.000 ;
    END
  END DA[9]
  PIN DB[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 174.800 4.510 176.800 ;
    END
  END DB[0]
  PIN DB[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 174.800 89.610 176.800 ;
    END
  END DB[10]
  PIN DB[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 174.800 98.350 176.800 ;
    END
  END DB[11]
  PIN DB[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 174.800 106.630 176.800 ;
    END
  END DB[12]
  PIN DB[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 174.800 115.370 176.800 ;
    END
  END DB[13]
  PIN DB[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 174.800 124.110 176.800 ;
    END
  END DB[14]
  PIN DB[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 174.800 132.390 176.800 ;
    END
  END DB[15]
  PIN DB[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 174.800 141.130 176.800 ;
    END
  END DB[16]
  PIN DB[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 174.800 149.410 176.800 ;
    END
  END DB[17]
  PIN DB[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 174.800 158.150 176.800 ;
    END
  END DB[18]
  PIN DB[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 174.800 166.430 176.800 ;
    END
  END DB[19]
  PIN DB[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 174.800 12.790 176.800 ;
    END
  END DB[1]
  PIN DB[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 174.800 175.170 176.800 ;
    END
  END DB[20]
  PIN DB[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 174.800 183.910 176.800 ;
    END
  END DB[21]
  PIN DB[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 174.800 192.190 176.800 ;
    END
  END DB[22]
  PIN DB[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 174.800 200.930 176.800 ;
    END
  END DB[23]
  PIN DB[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 174.800 209.210 176.800 ;
    END
  END DB[24]
  PIN DB[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 174.800 217.950 176.800 ;
    END
  END DB[25]
  PIN DB[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.950 174.800 226.230 176.800 ;
    END
  END DB[26]
  PIN DB[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 174.800 234.970 176.800 ;
    END
  END DB[27]
  PIN DB[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 174.800 243.710 176.800 ;
    END
  END DB[28]
  PIN DB[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 174.800 251.990 176.800 ;
    END
  END DB[29]
  PIN DB[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 174.800 21.530 176.800 ;
    END
  END DB[2]
  PIN DB[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 174.800 260.730 176.800 ;
    END
  END DB[30]
  PIN DB[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 174.800 269.010 176.800 ;
    END
  END DB[31]
  PIN DB[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 174.800 29.810 176.800 ;
    END
  END DB[3]
  PIN DB[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 174.800 38.550 176.800 ;
    END
  END DB[4]
  PIN DB[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 174.800 46.830 176.800 ;
    END
  END DB[5]
  PIN DB[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 174.800 55.570 176.800 ;
    END
  END DB[6]
  PIN DB[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 174.800 64.310 176.800 ;
    END
  END DB[7]
  PIN DB[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 174.800 72.590 176.800 ;
    END
  END DB[8]
  PIN DB[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 174.800 81.330 176.800 ;
    END
  END DB[9]
  PIN DW[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 0.000 164.130 2.000 ;
    END
  END DW[0]
  PIN DW[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 0.000 214.730 2.000 ;
    END
  END DW[10]
  PIN DW[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 0.000 219.790 2.000 ;
    END
  END DW[11]
  PIN DW[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 0.000 224.850 2.000 ;
    END
  END DW[12]
  PIN DW[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 0.000 229.910 2.000 ;
    END
  END DW[13]
  PIN DW[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 2.000 ;
    END
  END DW[14]
  PIN DW[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.750 0.000 240.030 2.000 ;
    END
  END DW[15]
  PIN DW[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 2.000 ;
    END
  END DW[16]
  PIN DW[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 0.000 250.150 2.000 ;
    END
  END DW[17]
  PIN DW[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 0.000 255.210 2.000 ;
    END
  END DW[18]
  PIN DW[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 0.000 260.270 2.000 ;
    END
  END DW[19]
  PIN DW[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 0.000 169.190 2.000 ;
    END
  END DW[1]
  PIN DW[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 0.000 265.330 2.000 ;
    END
  END DW[20]
  PIN DW[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 0.000 270.390 2.000 ;
    END
  END DW[21]
  PIN DW[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.170 0.000 275.450 2.000 ;
    END
  END DW[22]
  PIN DW[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 2.000 ;
    END
  END DW[23]
  PIN DW[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.290 0.000 285.570 2.000 ;
    END
  END DW[24]
  PIN DW[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.350 0.000 290.630 2.000 ;
    END
  END DW[25]
  PIN DW[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 0.000 295.690 2.000 ;
    END
  END DW[26]
  PIN DW[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.470 0.000 300.750 2.000 ;
    END
  END DW[27]
  PIN DW[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 0.000 305.810 2.000 ;
    END
  END DW[28]
  PIN DW[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.590 0.000 310.870 2.000 ;
    END
  END DW[29]
  PIN DW[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 2.000 ;
    END
  END DW[2]
  PIN DW[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 2.000 ;
    END
  END DW[30]
  PIN DW[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.710 0.000 320.990 2.000 ;
    END
  END DW[31]
  PIN DW[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.030 0.000 179.310 2.000 ;
    END
  END DW[3]
  PIN DW[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 2.000 ;
    END
  END DW[4]
  PIN DW[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 0.000 189.430 2.000 ;
    END
  END DW[5]
  PIN DW[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 0.000 194.490 2.000 ;
    END
  END DW[6]
  PIN DW[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.270 0.000 199.550 2.000 ;
    END
  END DW[7]
  PIN DW[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.330 0.000 204.610 2.000 ;
    END
  END DW[8]
  PIN DW[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 2.000 ;
    END
  END DW[9]
  PIN RA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.770 0.000 326.050 2.000 ;
    END
  END RA[0]
  PIN RA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 0.000 331.110 2.000 ;
    END
  END RA[1]
  PIN RA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 0.000 336.170 2.000 ;
    END
  END RA[2]
  PIN RA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.950 0.000 341.230 2.000 ;
    END
  END RA[3]
  PIN RA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.010 0.000 346.290 2.000 ;
    END
  END RA[4]
  PIN RB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 174.800 277.750 176.800 ;
    END
  END RB[0]
  PIN RB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 174.800 286.030 176.800 ;
    END
  END RB[1]
  PIN RB[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 174.800 294.770 176.800 ;
    END
  END RB[2]
  PIN RB[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.230 174.800 303.510 176.800 ;
    END
  END RB[3]
  PIN RB[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.510 174.800 311.790 176.800 ;
    END
  END RB[4]
  PIN RW[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.250 174.800 320.530 176.800 ;
    END
  END RW[0]
  PIN RW[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 174.800 328.810 176.800 ;
    END
  END RW[1]
  PIN RW[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 174.800 337.550 176.800 ;
    END
  END RW[2]
  PIN RW[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.550 174.800 345.830 176.800 ;
    END
  END RW[3]
  PIN RW[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 174.800 354.570 176.800 ;
    END
  END RW[4]
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 95.080 2.480 96.680 174.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 248.680 2.480 250.280 174.320 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.280 2.480 19.880 174.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.880 2.480 173.480 174.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.480 2.480 327.080 174.320 ;
    END
  END VPWR
  PIN WE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.130 0.000 356.410 2.000 ;
    END
  END WE
  OBS
      LAYER li1 ;
        RECT 2.760 2.635 356.040 174.165 ;
      LAYER met1 ;
        RECT 2.370 0.040 356.040 176.760 ;
      LAYER met2 ;
        RECT 2.390 174.520 3.950 176.790 ;
        RECT 4.790 174.520 12.230 176.790 ;
        RECT 13.070 174.520 20.970 176.790 ;
        RECT 21.810 174.520 29.250 176.790 ;
        RECT 30.090 174.520 37.990 176.790 ;
        RECT 38.830 174.520 46.270 176.790 ;
        RECT 47.110 174.520 55.010 176.790 ;
        RECT 55.850 174.520 63.750 176.790 ;
        RECT 64.590 174.520 72.030 176.790 ;
        RECT 72.870 174.520 80.770 176.790 ;
        RECT 81.610 174.520 89.050 176.790 ;
        RECT 89.890 174.520 97.790 176.790 ;
        RECT 98.630 174.520 106.070 176.790 ;
        RECT 106.910 174.520 114.810 176.790 ;
        RECT 115.650 174.520 123.550 176.790 ;
        RECT 124.390 174.520 131.830 176.790 ;
        RECT 132.670 174.520 140.570 176.790 ;
        RECT 141.410 174.520 148.850 176.790 ;
        RECT 149.690 174.520 157.590 176.790 ;
        RECT 158.430 174.520 165.870 176.790 ;
        RECT 166.710 174.520 174.610 176.790 ;
        RECT 175.450 174.520 183.350 176.790 ;
        RECT 184.190 174.520 191.630 176.790 ;
        RECT 192.470 174.520 200.370 176.790 ;
        RECT 201.210 174.520 208.650 176.790 ;
        RECT 209.490 174.520 217.390 176.790 ;
        RECT 218.230 174.520 225.670 176.790 ;
        RECT 226.510 174.520 234.410 176.790 ;
        RECT 235.250 174.520 243.150 176.790 ;
        RECT 243.990 174.520 251.430 176.790 ;
        RECT 252.270 174.520 260.170 176.790 ;
        RECT 261.010 174.520 268.450 176.790 ;
        RECT 269.290 174.520 277.190 176.790 ;
        RECT 278.030 174.520 285.470 176.790 ;
        RECT 286.310 174.520 294.210 176.790 ;
        RECT 295.050 174.520 302.950 176.790 ;
        RECT 303.790 174.520 311.230 176.790 ;
        RECT 312.070 174.520 319.970 176.790 ;
        RECT 320.810 174.520 328.250 176.790 ;
        RECT 329.090 174.520 336.990 176.790 ;
        RECT 337.830 174.520 345.270 176.790 ;
        RECT 346.110 174.520 354.010 176.790 ;
        RECT 354.850 174.520 356.410 176.790 ;
        RECT 2.390 2.280 356.410 174.520 ;
        RECT 2.950 0.010 6.710 2.280 ;
        RECT 7.550 0.010 11.770 2.280 ;
        RECT 12.610 0.010 16.830 2.280 ;
        RECT 17.670 0.010 21.890 2.280 ;
        RECT 22.730 0.010 26.950 2.280 ;
        RECT 27.790 0.010 32.010 2.280 ;
        RECT 32.850 0.010 37.070 2.280 ;
        RECT 37.910 0.010 42.130 2.280 ;
        RECT 42.970 0.010 47.190 2.280 ;
        RECT 48.030 0.010 52.250 2.280 ;
        RECT 53.090 0.010 57.310 2.280 ;
        RECT 58.150 0.010 62.370 2.280 ;
        RECT 63.210 0.010 67.430 2.280 ;
        RECT 68.270 0.010 72.490 2.280 ;
        RECT 73.330 0.010 77.550 2.280 ;
        RECT 78.390 0.010 82.610 2.280 ;
        RECT 83.450 0.010 87.670 2.280 ;
        RECT 88.510 0.010 92.730 2.280 ;
        RECT 93.570 0.010 97.790 2.280 ;
        RECT 98.630 0.010 102.850 2.280 ;
        RECT 103.690 0.010 107.910 2.280 ;
        RECT 108.750 0.010 112.970 2.280 ;
        RECT 113.810 0.010 118.030 2.280 ;
        RECT 118.870 0.010 123.090 2.280 ;
        RECT 123.930 0.010 128.150 2.280 ;
        RECT 128.990 0.010 133.210 2.280 ;
        RECT 134.050 0.010 138.270 2.280 ;
        RECT 139.110 0.010 143.330 2.280 ;
        RECT 144.170 0.010 148.390 2.280 ;
        RECT 149.230 0.010 153.450 2.280 ;
        RECT 154.290 0.010 158.510 2.280 ;
        RECT 159.350 0.010 163.570 2.280 ;
        RECT 164.410 0.010 168.630 2.280 ;
        RECT 169.470 0.010 173.690 2.280 ;
        RECT 174.530 0.010 178.750 2.280 ;
        RECT 179.590 0.010 183.810 2.280 ;
        RECT 184.650 0.010 188.870 2.280 ;
        RECT 189.710 0.010 193.930 2.280 ;
        RECT 194.770 0.010 198.990 2.280 ;
        RECT 199.830 0.010 204.050 2.280 ;
        RECT 204.890 0.010 209.110 2.280 ;
        RECT 209.950 0.010 214.170 2.280 ;
        RECT 215.010 0.010 219.230 2.280 ;
        RECT 220.070 0.010 224.290 2.280 ;
        RECT 225.130 0.010 229.350 2.280 ;
        RECT 230.190 0.010 234.410 2.280 ;
        RECT 235.250 0.010 239.470 2.280 ;
        RECT 240.310 0.010 244.530 2.280 ;
        RECT 245.370 0.010 249.590 2.280 ;
        RECT 250.430 0.010 254.650 2.280 ;
        RECT 255.490 0.010 259.710 2.280 ;
        RECT 260.550 0.010 264.770 2.280 ;
        RECT 265.610 0.010 269.830 2.280 ;
        RECT 270.670 0.010 274.890 2.280 ;
        RECT 275.730 0.010 279.950 2.280 ;
        RECT 280.790 0.010 285.010 2.280 ;
        RECT 285.850 0.010 290.070 2.280 ;
        RECT 290.910 0.010 295.130 2.280 ;
        RECT 295.970 0.010 300.190 2.280 ;
        RECT 301.030 0.010 305.250 2.280 ;
        RECT 306.090 0.010 310.310 2.280 ;
        RECT 311.150 0.010 315.370 2.280 ;
        RECT 316.210 0.010 320.430 2.280 ;
        RECT 321.270 0.010 325.490 2.280 ;
        RECT 326.330 0.010 330.550 2.280 ;
        RECT 331.390 0.010 335.610 2.280 ;
        RECT 336.450 0.010 340.670 2.280 ;
        RECT 341.510 0.010 345.730 2.280 ;
        RECT 346.570 0.010 350.790 2.280 ;
        RECT 351.630 0.010 355.850 2.280 ;
      LAYER met3 ;
        RECT 2.365 0.175 356.435 176.625 ;
      LAYER met4 ;
        RECT 98.735 174.720 342.865 176.625 ;
        RECT 98.735 2.080 171.480 174.720 ;
        RECT 173.880 2.080 248.280 174.720 ;
        RECT 250.680 2.080 325.080 174.720 ;
        RECT 327.480 2.080 342.865 174.720 ;
        RECT 98.735 1.535 342.865 2.080 ;
  END
END DFFRF_2R1W
END LIBRARY

